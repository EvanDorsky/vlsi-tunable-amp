magic
tech scmos
timestamp 1417990464
<< ntransistor >>
rect 0 24 4 26
<< ptransistor >>
rect 0 0 4 2
<< ndiffusion >>
rect 0 26 4 27
rect 0 23 4 24
<< pdiffusion >>
rect 0 2 4 3
rect 0 -1 4 0
<< ndcontact >>
rect 0 27 4 31
rect 0 19 4 23
<< pdcontact >>
rect 0 3 4 7
rect 0 -5 4 -1
<< polysilicon >>
rect -3 24 0 26
rect 4 24 6 26
rect -3 2 -1 24
rect -3 0 0 2
rect 4 0 6 2
<< metal1 >>
rect -3 27 0 31
rect 4 27 6 31
rect 0 15 4 19
rect 0 11 6 15
rect 0 7 4 11
rect -3 -5 0 -1
rect 4 -5 6 -1
<< labels >>
rlabel polysilicon -3 12 -2 14 3 A
rlabel metal1 5 11 6 15 7 Z
rlabel metal1 -3 -5 -2 -1 2 Gnd
rlabel metal1 -3 27 -2 31 4 Vdd
<< end >>
