magic
tech scmos
magscale 1 3
timestamp 1419146600
<< metal1 >>
rect 2074 7175 2104 7185
rect 2034 7165 2134 7175
rect 1994 7155 2154 7165
rect 1974 7145 2174 7155
rect 1954 7135 2184 7145
rect 1934 7125 2194 7135
rect 1924 7115 2304 7125
rect 1924 7105 2314 7115
rect 1934 7095 2334 7105
rect 1934 7085 2344 7095
rect 1804 7075 1824 7085
rect 1934 7075 2364 7085
rect 1794 7065 1844 7075
rect 1934 7065 2394 7075
rect 1644 7055 1674 7065
rect 1634 7045 1674 7055
rect 1794 7045 1864 7065
rect 1934 7055 2414 7065
rect 1924 7045 2424 7055
rect 1624 7035 1664 7045
rect 1604 7025 1664 7035
rect 1804 7035 1864 7045
rect 1914 7035 2434 7045
rect 2544 7035 2574 7045
rect 1804 7025 1874 7035
rect 1904 7025 2464 7035
rect 2524 7025 2614 7035
rect 2674 7025 2744 7035
rect 1594 7015 1664 7025
rect 1814 7015 2754 7025
rect 1574 7005 1714 7015
rect 1814 7005 2764 7015
rect 1554 6995 1714 7005
rect 1524 6985 1714 6995
rect 1504 6975 1714 6985
rect 1494 6965 1714 6975
rect 1844 6995 2804 7005
rect 2904 6995 3014 7005
rect 1844 6985 2814 6995
rect 2884 6985 3024 6995
rect 1844 6975 2834 6985
rect 2844 6975 3014 6985
rect 1844 6965 3014 6975
rect 1504 6945 1704 6965
rect 1824 6955 3004 6965
rect 1804 6945 3004 6955
rect 3264 6945 3304 6955
rect 1444 6935 1454 6945
rect 1434 6925 1454 6935
rect 1424 6905 1454 6925
rect 1514 6935 1704 6945
rect 1794 6935 3004 6945
rect 3254 6935 3314 6945
rect 1514 6925 1744 6935
rect 1774 6925 3004 6935
rect 1514 6915 3004 6925
rect 1514 6905 3014 6915
rect 3104 6905 3114 6915
rect 1414 6885 1444 6905
rect 1504 6895 1664 6905
rect 1674 6895 3224 6905
rect 1494 6885 1634 6895
rect 1694 6885 3234 6895
rect 1404 6875 1444 6885
rect 1484 6875 1634 6885
rect 1414 6865 1444 6875
rect 1474 6865 1644 6875
rect 1704 6865 3244 6885
rect 1404 6855 1654 6865
rect 1694 6855 2954 6865
rect 2964 6855 3254 6865
rect 1374 6845 2944 6855
rect 1344 6835 2944 6845
rect 2964 6835 3264 6855
rect 1304 6825 2874 6835
rect 2964 6825 3274 6835
rect 1304 6815 2854 6825
rect 2954 6815 3274 6825
rect 1294 6805 2854 6815
rect 2944 6805 3274 6815
rect 1284 6795 2874 6805
rect 2934 6795 3284 6805
rect 3464 6795 3514 6805
rect 1284 6785 2534 6795
rect 2574 6785 3284 6795
rect 3424 6785 3524 6795
rect 1274 6775 2524 6785
rect 1264 6765 2514 6775
rect 2574 6765 3294 6785
rect 3404 6775 3534 6785
rect 3404 6765 3544 6775
rect 1204 6755 2114 6765
rect 2124 6755 2334 6765
rect 2344 6755 2504 6765
rect 1184 6735 2104 6755
rect 2124 6745 2314 6755
rect 2354 6745 2504 6755
rect 2574 6745 3304 6765
rect 3394 6755 3564 6765
rect 3394 6745 3574 6755
rect 2124 6735 2304 6745
rect 2344 6735 2504 6745
rect 2564 6735 3324 6745
rect 3394 6735 3584 6745
rect 1174 6725 2104 6735
rect 2134 6725 2304 6735
rect 2334 6725 3334 6735
rect 3394 6725 3594 6735
rect 1174 6715 2114 6725
rect 2124 6715 2294 6725
rect 2324 6715 3344 6725
rect 3394 6715 3604 6725
rect 1174 6705 2154 6715
rect 2194 6705 2294 6715
rect 2314 6705 3354 6715
rect 3394 6705 3614 6715
rect 1174 6695 2144 6705
rect 2194 6695 2284 6705
rect 2304 6695 3364 6705
rect 3384 6695 3614 6705
rect 1174 6675 2134 6695
rect 2194 6685 2274 6695
rect 2184 6675 2274 6685
rect 2304 6685 2514 6695
rect 2544 6685 3624 6695
rect 1164 6665 2124 6675
rect 2174 6665 2264 6675
rect 1164 6655 2104 6665
rect 2174 6655 2244 6665
rect 2304 6655 2504 6685
rect 2554 6665 3634 6685
rect 2554 6655 3644 6665
rect 1144 6645 2084 6655
rect 2174 6645 2224 6655
rect 1134 6635 2074 6645
rect 1124 6625 1994 6635
rect 2044 6625 2064 6635
rect 2174 6625 2214 6645
rect 2294 6635 2504 6655
rect 2544 6645 3634 6655
rect 2544 6635 3254 6645
rect 3284 6635 3644 6645
rect 3674 6635 3684 6645
rect 2284 6625 2514 6635
rect 2534 6625 3254 6635
rect 3304 6625 3694 6635
rect 1104 6615 1954 6625
rect 2164 6615 2214 6625
rect 2274 6615 3244 6625
rect 1104 6605 1934 6615
rect 2154 6605 2224 6615
rect 2264 6605 2784 6615
rect 2814 6605 3244 6615
rect 3314 6615 3694 6625
rect 3314 6605 3534 6615
rect 3564 6605 3694 6615
rect 1094 6595 1924 6605
rect 2054 6595 2064 6605
rect 2144 6595 2774 6605
rect 2814 6595 3254 6605
rect 3294 6595 3524 6605
rect 3574 6595 3684 6605
rect 1084 6585 1924 6595
rect 2044 6585 2074 6595
rect 2134 6585 2764 6595
rect 2804 6585 3254 6595
rect 3274 6585 3454 6595
rect 1074 6575 1934 6585
rect 2034 6575 2084 6585
rect 2114 6575 2754 6585
rect 2794 6575 3454 6585
rect 3464 6585 3504 6595
rect 3614 6585 3664 6595
rect 3464 6575 3494 6585
rect 1074 6565 1984 6575
rect 2024 6565 2744 6575
rect 2774 6565 3494 6575
rect 1074 6555 2734 6565
rect 2754 6555 3484 6565
rect 1074 6535 2474 6555
rect 2494 6545 2724 6555
rect 2744 6545 3494 6555
rect 2504 6535 3494 6545
rect 1074 6525 2464 6535
rect 1084 6505 2464 6525
rect 2504 6515 3504 6535
rect 2494 6505 3504 6515
rect 3654 6525 3684 6535
rect 3654 6505 3694 6525
rect 1084 6495 1524 6505
rect 1554 6495 3514 6505
rect 3654 6495 3704 6505
rect 1084 6485 1514 6495
rect 1564 6485 1914 6495
rect 1934 6485 3514 6495
rect 3644 6485 3704 6495
rect 1084 6475 1444 6485
rect 1494 6475 1504 6485
rect 1564 6475 1904 6485
rect 1934 6475 3524 6485
rect 1084 6465 1434 6475
rect 1084 6435 1424 6465
rect 1464 6445 1504 6455
rect 1574 6445 1894 6475
rect 1934 6465 2334 6475
rect 2344 6465 3534 6475
rect 3634 6465 3704 6485
rect 1924 6445 2334 6465
rect 2354 6445 3554 6465
rect 3644 6445 3704 6465
rect 1434 6435 1514 6445
rect 1094 6425 1514 6435
rect 1584 6435 1904 6445
rect 1914 6435 2634 6445
rect 1584 6425 2634 6435
rect 2664 6425 3564 6445
rect 3634 6425 3704 6445
rect 1104 6405 1524 6425
rect 1584 6415 1834 6425
rect 1874 6415 2634 6425
rect 2654 6415 3564 6425
rect 3614 6415 3704 6425
rect 1104 6395 1384 6405
rect 1424 6395 1524 6405
rect 1574 6395 1834 6415
rect 1864 6405 3564 6415
rect 3604 6405 3704 6415
rect 1854 6395 3684 6405
rect 1104 6385 1364 6395
rect 1434 6385 1524 6395
rect 1094 6375 1354 6385
rect 1424 6375 1534 6385
rect 1564 6375 3674 6395
rect 3684 6375 3714 6385
rect 3804 6375 3864 6385
rect 1094 6365 1344 6375
rect 1414 6365 3724 6375
rect 3794 6365 3874 6375
rect 1094 6355 1334 6365
rect 1404 6355 3744 6365
rect 3784 6355 3874 6365
rect 1084 6345 1574 6355
rect 1614 6345 3874 6355
rect 1084 6335 1554 6345
rect 1074 6325 1444 6335
rect 1494 6325 1544 6335
rect 1624 6325 3874 6345
rect 1064 6315 1434 6325
rect 1054 6305 1424 6315
rect 1614 6305 3874 6325
rect 984 6295 1004 6305
rect 1044 6295 1414 6305
rect 1604 6295 3874 6305
rect 954 6285 1404 6295
rect 944 6275 1394 6285
rect 1604 6275 3864 6295
rect 934 6265 1384 6275
rect 1594 6265 3864 6275
rect 924 6255 1384 6265
rect 1484 6255 1504 6265
rect 1574 6255 2484 6265
rect 2524 6255 2654 6265
rect 2704 6255 3874 6265
rect 904 6245 1394 6255
rect 1404 6245 1514 6255
rect 1564 6245 2474 6255
rect 2534 6245 2624 6255
rect 894 6235 2474 6245
rect 2544 6235 2624 6245
rect 874 6225 2474 6235
rect 864 6215 2474 6225
rect 2554 6215 2624 6235
rect 2714 6245 3884 6255
rect 2714 6235 3704 6245
rect 3714 6235 3884 6245
rect 2714 6225 3684 6235
rect 3724 6225 3894 6235
rect 2704 6215 3684 6225
rect 854 6205 2484 6215
rect 2554 6205 2604 6215
rect 2684 6205 3684 6215
rect 3734 6205 3894 6225
rect 764 6195 794 6205
rect 854 6195 2594 6205
rect 2674 6195 3684 6205
rect 754 6185 804 6195
rect 744 6175 804 6185
rect 854 6185 2584 6195
rect 744 6165 794 6175
rect 734 6145 794 6165
rect 854 6165 2594 6185
rect 2664 6175 3684 6195
rect 2664 6165 3264 6175
rect 3274 6165 3694 6175
rect 854 6155 2604 6165
rect 2664 6155 3694 6165
rect 844 6145 2614 6155
rect 2654 6145 3694 6155
rect 3724 6145 3894 6205
rect 734 6135 774 6145
rect 834 6135 3694 6145
rect 734 6125 764 6135
rect 824 6115 3704 6135
rect 3734 6125 3894 6145
rect 814 6105 2404 6115
rect 2414 6105 3704 6115
rect 814 6095 2374 6105
rect 2434 6095 3704 6105
rect 814 6085 2354 6095
rect 2444 6085 3704 6095
rect 804 6075 2344 6085
rect 2454 6075 3704 6085
rect 804 6055 2334 6075
rect 804 6045 2324 6055
rect 804 6025 2334 6045
rect 794 6015 2334 6025
rect 2444 6035 3704 6075
rect 3744 6095 3894 6125
rect 3744 6075 3884 6095
rect 3744 6065 3874 6075
rect 3754 6055 3814 6065
rect 3764 6045 3804 6055
rect 3784 6035 3794 6045
rect 2444 6025 2854 6035
rect 2894 6025 3694 6035
rect 2444 6015 2844 6025
rect 2934 6015 3694 6025
rect 784 6005 2334 6015
rect 724 5995 2334 6005
rect 2454 5995 2834 6015
rect 2964 6005 3694 6015
rect 2984 5995 3684 6005
rect 714 5975 2344 5995
rect 2454 5985 2824 5995
rect 2994 5985 3684 5995
rect 714 5965 2354 5975
rect 2464 5965 2824 5985
rect 2974 5975 3784 5985
rect 2934 5965 3854 5975
rect 704 5955 2354 5965
rect 704 5945 2344 5955
rect 2454 5945 2814 5965
rect 2884 5955 3904 5965
rect 3994 5955 4024 5965
rect 2854 5945 4024 5955
rect 704 5935 2334 5945
rect 2504 5935 2814 5945
rect 2824 5935 4024 5945
rect 704 5925 2324 5935
rect 2514 5925 4014 5935
rect 704 5915 2314 5925
rect 2524 5915 4014 5925
rect 704 5905 2304 5915
rect 2534 5905 4004 5915
rect 694 5885 2294 5905
rect 2554 5895 2594 5905
rect 2674 5895 3994 5905
rect 2694 5885 3984 5895
rect 694 5875 2284 5885
rect 2674 5875 3964 5885
rect 684 5865 2274 5875
rect 2654 5865 3934 5875
rect 684 5855 2264 5865
rect 2634 5855 3884 5865
rect 694 5845 2214 5855
rect 2614 5845 3864 5855
rect 694 5835 2184 5845
rect 2594 5835 3854 5845
rect 704 5825 2134 5835
rect 2574 5825 3844 5835
rect 704 5815 2114 5825
rect 2564 5815 3834 5825
rect 704 5805 2104 5815
rect 2544 5805 3834 5815
rect 704 5795 2084 5805
rect 2534 5795 2764 5805
rect 2794 5795 3824 5805
rect 694 5785 2064 5795
rect 2514 5785 2754 5795
rect 2804 5785 3824 5795
rect 694 5765 2044 5785
rect 2504 5775 2744 5785
rect 2824 5775 3814 5785
rect 2524 5765 2724 5775
rect 2834 5765 3664 5775
rect 3704 5765 3814 5775
rect 694 5755 2034 5765
rect 2534 5755 2664 5765
rect 2844 5755 3644 5765
rect 3734 5755 3814 5765
rect 694 5745 2024 5755
rect 2544 5745 2614 5755
rect 2954 5745 3244 5755
rect 3304 5745 3614 5755
rect 3754 5745 3814 5755
rect 684 5715 2024 5745
rect 2554 5735 2594 5745
rect 2964 5735 3234 5745
rect 3324 5735 3524 5745
rect 2974 5725 3214 5735
rect 3344 5725 3494 5735
rect 2984 5715 3194 5725
rect 3364 5715 3464 5725
rect 3764 5715 3814 5745
rect 674 5705 2024 5715
rect 664 5695 774 5705
rect 824 5695 2024 5705
rect 3004 5705 3174 5715
rect 3384 5705 3444 5715
rect 3004 5695 3124 5705
rect 3774 5695 3824 5715
rect 654 5685 714 5695
rect 734 5685 744 5695
rect 654 5675 674 5685
rect 894 5675 2024 5695
rect 3014 5685 3104 5695
rect 3774 5685 3834 5695
rect 2384 5675 2424 5685
rect 3024 5675 3084 5685
rect 3784 5675 3834 5685
rect 654 5665 664 5675
rect 894 5665 2034 5675
rect 2374 5665 2424 5675
rect 894 5655 2044 5665
rect 2374 5655 2434 5665
rect 3784 5655 3844 5675
rect 894 5645 2054 5655
rect 884 5635 2064 5645
rect 2374 5635 2424 5655
rect 3794 5645 3844 5655
rect 884 5625 2074 5635
rect 2374 5625 2414 5635
rect 3794 5625 3834 5645
rect 874 5615 2084 5625
rect 864 5605 2094 5615
rect 854 5595 2094 5605
rect 854 5585 2104 5595
rect 844 5575 2104 5585
rect 844 5565 2114 5575
rect 834 5555 2114 5565
rect 2264 5555 2284 5565
rect 824 5535 2124 5555
rect 2254 5545 2284 5555
rect 2244 5535 2284 5545
rect 814 5525 1964 5535
rect 1984 5525 2134 5535
rect 2234 5525 2284 5535
rect 814 5505 1954 5525
rect 1994 5515 2134 5525
rect 2224 5515 2274 5525
rect 1984 5505 2134 5515
rect 2214 5505 2274 5515
rect 804 5485 2144 5505
rect 2204 5495 2274 5505
rect 2194 5485 2274 5495
rect 804 5475 2174 5485
rect 2184 5475 2274 5485
rect 794 5455 2284 5475
rect 784 5445 2154 5455
rect 2164 5445 2294 5455
rect 774 5425 2294 5445
rect 4094 5435 4144 5445
rect 4044 5425 4174 5435
rect 764 5405 2294 5425
rect 3804 5415 3874 5425
rect 4004 5415 4184 5425
rect 3784 5405 4184 5415
rect 754 5375 2294 5405
rect 3764 5395 4184 5405
rect 3754 5385 4184 5395
rect 3734 5375 4184 5385
rect 754 5355 2304 5375
rect 3714 5365 4184 5375
rect 3704 5355 4184 5365
rect 754 5345 2314 5355
rect 3684 5345 4184 5355
rect 764 5335 2324 5345
rect 3664 5335 4184 5345
rect 764 5325 2334 5335
rect 3654 5325 4184 5335
rect 774 5315 2344 5325
rect 3634 5315 4184 5325
rect 774 5305 2354 5315
rect 3614 5305 4174 5315
rect 804 5295 2364 5305
rect 3594 5295 4174 5305
rect 814 5285 2364 5295
rect 3574 5285 4044 5295
rect 4064 5285 4164 5295
rect 824 5275 2374 5285
rect 3554 5275 4034 5285
rect 4074 5275 4164 5285
rect 834 5255 2374 5275
rect 3154 5265 3264 5275
rect 3314 5265 3354 5275
rect 3534 5265 4034 5275
rect 3134 5255 3414 5265
rect 3514 5255 4034 5265
rect 844 5245 2374 5255
rect 3094 5245 3464 5255
rect 3494 5245 4034 5255
rect 844 5225 2364 5245
rect 3074 5235 4034 5245
rect 3054 5225 4034 5235
rect 4084 5225 4154 5275
rect 844 5195 2354 5225
rect 3014 5215 4024 5225
rect 3004 5205 4024 5215
rect 4094 5205 4154 5225
rect 2984 5195 4014 5205
rect 854 5185 2364 5195
rect 2964 5185 4014 5195
rect 854 5175 2374 5185
rect 2944 5175 4014 5185
rect 864 5165 2444 5175
rect 2934 5165 4014 5175
rect 864 5155 2514 5165
rect 2914 5155 4014 5165
rect 874 5145 2534 5155
rect 2604 5154 2634 5155
rect 2595 5145 2634 5154
rect 2884 5145 4014 5155
rect 884 5135 2604 5145
rect 2874 5135 4014 5145
rect 884 5125 2564 5135
rect 2854 5125 4014 5135
rect 884 5115 2514 5125
rect 2844 5115 4014 5125
rect 884 5105 2484 5115
rect 2824 5105 4014 5115
rect 884 5095 2464 5105
rect 2814 5095 4014 5105
rect 4084 5105 4154 5205
rect 4084 5095 4144 5105
rect 884 5085 2454 5095
rect 2794 5085 4014 5095
rect 884 5075 2424 5085
rect 2794 5075 4024 5085
rect 884 5065 2404 5075
rect 2774 5065 4024 5075
rect 894 5055 2404 5065
rect 894 5015 2414 5055
rect 2764 5045 4024 5065
rect 4074 5055 4144 5095
rect 2754 5035 3514 5045
rect 3534 5035 4024 5045
rect 2744 5025 3504 5035
rect 3554 5025 4024 5035
rect 4084 5035 4144 5055
rect 4084 5025 4134 5035
rect 2744 5015 3494 5025
rect 3574 5015 4024 5025
rect 4074 5015 4134 5025
rect 904 5005 2414 5015
rect 2534 5005 2584 5015
rect 2694 5005 2714 5015
rect 904 4995 2424 5005
rect 2524 4995 2624 5005
rect 2674 4995 2714 5005
rect 2734 5005 3494 5015
rect 3584 5005 4024 5015
rect 2734 4995 3484 5005
rect 904 4985 2714 4995
rect 2724 4985 3484 4995
rect 3594 4985 4024 5005
rect 4084 4995 4134 5015
rect 4074 4985 4124 4995
rect 914 4975 1404 4985
rect 1454 4975 3484 4985
rect 3614 4975 4024 4985
rect 924 4965 1374 4975
rect 1474 4965 3474 4975
rect 3624 4965 4014 4975
rect 4054 4965 4124 4985
rect 924 4955 1364 4965
rect 1484 4955 3474 4965
rect 934 4945 1354 4955
rect 1494 4945 3474 4955
rect 3634 4955 4024 4965
rect 4054 4955 4114 4965
rect 3634 4945 4114 4955
rect 934 4935 1344 4945
rect 1504 4935 3474 4945
rect 3644 4935 4114 4945
rect 944 4915 1334 4935
rect 1514 4925 3474 4935
rect 1524 4915 3474 4925
rect 3654 4915 4104 4935
rect 954 4905 1324 4915
rect 1544 4905 3474 4915
rect 954 4895 1314 4905
rect 1554 4895 3474 4905
rect 3664 4895 4094 4915
rect 954 4875 1304 4895
rect 1584 4885 3464 4895
rect 3674 4885 4094 4895
rect 1604 4875 3464 4885
rect 964 4855 1304 4875
rect 1624 4865 3464 4875
rect 3684 4865 4084 4885
rect 1634 4855 3464 4865
rect 3694 4855 4074 4865
rect 964 4835 1294 4855
rect 1644 4845 3454 4855
rect 1654 4835 3454 4845
rect 3704 4845 4074 4855
rect 3704 4835 4064 4845
rect 974 4815 1294 4835
rect 1674 4815 3454 4835
rect 3714 4825 4054 4835
rect 984 4805 1294 4815
rect 1684 4805 3444 4815
rect 3724 4805 4044 4825
rect 984 4795 1304 4805
rect 994 4775 1304 4795
rect 1004 4735 1304 4775
rect 1684 4795 2294 4805
rect 2434 4795 3444 4805
rect 3734 4795 4034 4805
rect 1684 4785 2244 4795
rect 2494 4785 3444 4795
rect 3744 4785 4024 4795
rect 1684 4775 2174 4785
rect 2514 4775 2554 4785
rect 2594 4775 3434 4785
rect 3744 4775 4014 4785
rect 1684 4755 2154 4775
rect 2614 4765 3434 4775
rect 3754 4765 4004 4775
rect 2624 4755 3434 4765
rect 3764 4755 3994 4765
rect 1684 4735 2144 4755
rect 2634 4735 3424 4755
rect 3774 4745 3974 4755
rect 3784 4735 3954 4745
rect 1004 4715 1314 4735
rect 1674 4725 2144 4735
rect 994 4705 1314 4715
rect 1664 4715 1744 4725
rect 1764 4715 2154 4725
rect 2644 4715 3424 4735
rect 3794 4725 3934 4735
rect 3814 4715 3914 4725
rect 1664 4705 1714 4715
rect 994 4685 1324 4705
rect 1674 4695 1704 4705
rect 1794 4695 2164 4715
rect 2654 4695 3424 4715
rect 3824 4705 3894 4715
rect 3844 4695 3884 4705
rect 1784 4685 2174 4695
rect 2654 4685 3414 4695
rect 994 4675 1334 4685
rect 984 4665 1334 4675
rect 1784 4675 2184 4685
rect 1784 4665 2194 4675
rect 2664 4665 3414 4685
rect 984 4655 1344 4665
rect 1784 4655 2204 4665
rect 2664 4655 3404 4665
rect 984 4635 1354 4655
rect 1774 4645 2224 4655
rect 2674 4645 3404 4655
rect 1774 4635 1804 4645
rect 1854 4635 2234 4645
rect 2674 4635 3394 4645
rect 984 4615 1364 4635
rect 1774 4625 1794 4635
rect 1874 4625 2234 4635
rect 1774 4615 1784 4625
rect 1894 4615 2234 4625
rect 984 4605 1374 4615
rect 1914 4605 2234 4615
rect 2684 4605 3374 4635
rect 994 4585 1384 4605
rect 994 4575 1394 4585
rect 1924 4575 2234 4605
rect 2694 4595 3364 4605
rect 2704 4585 3364 4595
rect 2714 4575 3364 4585
rect 1004 4565 1394 4575
rect 1014 4555 1404 4565
rect 1764 4555 1774 4575
rect 1934 4555 2234 4575
rect 2724 4565 3354 4575
rect 2744 4555 3254 4565
rect 3284 4555 3354 4565
rect 1024 4545 1414 4555
rect 1764 4545 1784 4555
rect 1044 4535 1464 4545
rect 1064 4525 1464 4535
rect 1764 4525 1794 4545
rect 1934 4535 2244 4555
rect 2744 4545 3234 4555
rect 3294 4545 3354 4555
rect 2764 4535 3194 4545
rect 3304 4535 3354 4545
rect 1934 4525 2254 4535
rect 2774 4525 3164 4535
rect 3304 4525 3364 4535
rect 1074 4515 1474 4525
rect 1764 4515 1804 4525
rect 1074 4505 1484 4515
rect 1764 4505 1814 4515
rect 1944 4505 2254 4525
rect 2844 4515 3144 4525
rect 2924 4505 3124 4515
rect 3314 4505 3364 4525
rect 3514 4515 3634 4525
rect 3494 4505 3654 4515
rect 1084 4495 1494 4505
rect 1774 4495 1844 4505
rect 1144 4485 1504 4495
rect 1784 4485 1854 4495
rect 1944 4485 2244 4505
rect 2944 4495 3094 4505
rect 3314 4495 3374 4505
rect 3484 4495 3674 4505
rect 2974 4485 3054 4495
rect 3324 4485 3404 4495
rect 3464 4485 3684 4495
rect 1174 4475 1514 4485
rect 1784 4475 1874 4485
rect 1944 4475 2234 4485
rect 2294 4475 2354 4485
rect 3324 4475 3424 4485
rect 3434 4475 3694 4485
rect 1194 4465 1514 4475
rect 1214 4455 1524 4465
rect 1794 4455 1884 4475
rect 1214 4445 1534 4455
rect 1814 4445 1874 4455
rect 1944 4445 2224 4475
rect 2294 4445 2364 4475
rect 3334 4465 3694 4475
rect 3344 4455 3694 4465
rect 3364 4445 3694 4455
rect 1224 4435 1544 4445
rect 1944 4435 2234 4445
rect 2294 4435 2354 4445
rect 3384 4435 3694 4445
rect 1224 4425 1554 4435
rect 1214 4415 1554 4425
rect 1934 4415 2234 4435
rect 2284 4425 2344 4435
rect 3404 4425 3684 4435
rect 2284 4415 2334 4425
rect 3414 4415 3534 4425
rect 3604 4415 3684 4425
rect 1214 4405 1564 4415
rect 1214 4385 1574 4405
rect 1924 4395 2234 4415
rect 2274 4405 2334 4415
rect 2274 4395 2314 4405
rect 3614 4395 3684 4415
rect 1214 4375 1584 4385
rect 1914 4375 2244 4395
rect 3614 4385 3674 4395
rect 3614 4375 3664 4385
rect 1214 4365 1594 4375
rect 1924 4365 2254 4375
rect 1224 4355 1604 4365
rect 1934 4355 2254 4365
rect 1224 4345 1614 4355
rect 1944 4345 2254 4355
rect 1224 4335 1624 4345
rect 1954 4335 2264 4345
rect 2314 4335 2334 4345
rect 1234 4325 1634 4335
rect 1954 4325 2274 4335
rect 2304 4325 2334 4335
rect 1234 4315 1654 4325
rect 1964 4315 2284 4325
rect 2294 4315 2334 4325
rect 1254 4305 1664 4315
rect 1964 4305 2314 4315
rect 1264 4295 1684 4305
rect 1284 4285 1694 4295
rect 1314 4275 1704 4285
rect 1324 4265 1714 4275
rect 1974 4265 2304 4305
rect 1324 4255 1724 4265
rect 1964 4255 2304 4265
rect 1314 4245 1744 4255
rect 1954 4245 2304 4255
rect 3824 4245 3844 4255
rect 1304 4235 1764 4245
rect 1934 4235 2364 4245
rect 3784 4235 3844 4245
rect 1304 4225 1794 4235
rect 1914 4225 2374 4235
rect 3764 4225 3844 4235
rect 1304 4215 1834 4225
rect 1894 4215 2374 4225
rect 1304 4205 2374 4215
rect 3744 4205 3844 4225
rect 1314 4195 2374 4205
rect 3454 4195 3504 4205
rect 3674 4195 3844 4205
rect 1314 4185 2384 4195
rect 3414 4185 3524 4195
rect 3574 4185 3834 4195
rect 1324 4175 2384 4185
rect 3364 4175 3754 4185
rect 1324 4165 2324 4175
rect 2334 4165 2384 4175
rect 3314 4165 3734 4175
rect 1334 4155 2324 4165
rect 1344 4145 2324 4155
rect 2354 4145 2374 4165
rect 3224 4155 3684 4165
rect 3204 4145 3464 4155
rect 3494 4145 3674 4155
rect 1354 4135 2334 4145
rect 1364 4125 2334 4135
rect 3194 4135 3424 4145
rect 3194 4125 3394 4135
rect 1364 4115 2344 4125
rect 3184 4115 3384 4125
rect 1374 4105 2354 4115
rect 1394 4095 2354 4105
rect 3184 4105 3344 4115
rect 3184 4095 3304 4105
rect 1404 4085 2364 4095
rect 1424 4075 2374 4085
rect 1434 4065 2384 4075
rect 1444 4055 2394 4065
rect 1454 4045 2404 4055
rect 1464 4035 2414 4045
rect 1474 4025 2414 4035
rect 3664 4025 3734 4035
rect 1484 4015 2424 4025
rect 3624 4015 3734 4025
rect 1494 4005 2434 4015
rect 3574 4005 3744 4015
rect 1514 3995 2444 4005
rect 3504 3995 3734 4005
rect 1554 3985 2454 3995
rect 3484 3985 3734 3995
rect 1574 3975 1614 3985
rect 1654 3975 2464 3985
rect 3464 3975 3724 3985
rect 1664 3965 2464 3975
rect 3434 3965 3714 3975
rect 1664 3955 2474 3965
rect 3424 3955 3694 3965
rect 1674 3945 2484 3955
rect 3434 3945 3664 3955
rect 1674 3935 2504 3945
rect 3464 3935 3504 3945
rect 1684 3925 2524 3935
rect 1704 3915 2574 3925
rect 1734 3905 2584 3915
rect 1784 3895 2594 3905
rect 1804 3885 2614 3895
rect 1804 3875 2634 3885
rect 1804 3865 2654 3875
rect 1804 3855 2684 3865
rect 1804 3845 2734 3855
rect 1804 3835 2754 3845
rect 1804 3825 2804 3835
rect 1804 3815 2864 3825
rect 1804 3805 2884 3815
rect 1804 3795 2894 3805
rect 1804 3785 2934 3795
rect 1804 3765 2944 3785
rect 3344 3765 3404 3775
rect 1804 3755 2954 3765
rect 3324 3755 3394 3765
rect 1804 3745 2964 3755
rect 3024 3745 3034 3755
rect 3294 3745 3384 3755
rect 1804 3735 2974 3745
rect 2994 3735 3084 3745
rect 3104 3735 3144 3745
rect 3214 3735 3374 3745
rect 1804 3725 3364 3735
rect 1804 3715 3344 3725
rect 1804 3705 3334 3715
rect 1794 3695 3314 3705
rect 1794 3685 3294 3695
rect 1794 3675 3284 3685
rect 1794 3665 3274 3675
rect 1794 3655 3264 3665
rect 1794 3645 3254 3655
rect 1794 3635 3244 3645
rect 3824 3635 3844 3645
rect 1794 3625 3234 3635
rect 3794 3625 3854 3635
rect 1784 3615 3234 3625
rect 3774 3615 3834 3625
rect 1784 3605 3224 3615
rect 3764 3605 3824 3615
rect 1784 3595 3214 3605
rect 3754 3595 3814 3605
rect 1774 3585 3204 3595
rect 3764 3585 3794 3595
rect 1774 3575 3194 3585
rect 1774 3565 3184 3575
rect 1764 3555 3184 3565
rect 1764 3545 2174 3555
rect 2184 3545 3174 3555
rect 1754 3535 2164 3545
rect 2194 3535 3164 3545
rect 1744 3525 2164 3535
rect 2264 3525 3154 3535
rect 1744 3515 2154 3525
rect 2274 3515 3144 3525
rect 1734 3505 2154 3515
rect 2284 3505 3134 3515
rect 1734 3495 2144 3505
rect 2304 3495 3124 3505
rect 1724 3485 2144 3495
rect 2324 3485 3114 3495
rect 1724 3475 2114 3485
rect 2344 3475 3104 3485
rect 1714 3465 2104 3475
rect 2354 3465 3094 3475
rect 1704 3455 2094 3465
rect 2374 3455 3084 3465
rect 1694 3435 2094 3455
rect 2384 3445 3074 3455
rect 2394 3435 3054 3445
rect 1684 3425 2094 3435
rect 2404 3425 3044 3435
rect 1454 3415 1524 3425
rect 1694 3415 1714 3425
rect 1764 3415 2104 3425
rect 2404 3415 3034 3425
rect 1434 3405 1554 3415
rect 1764 3405 2144 3415
rect 2404 3405 3014 3415
rect 1414 3395 1564 3405
rect 1774 3395 2154 3405
rect 2414 3395 3004 3405
rect 1404 3385 1554 3395
rect 1814 3385 2144 3395
rect 2424 3385 2994 3395
rect 1384 3375 1554 3385
rect 1854 3375 2114 3385
rect 2454 3375 2984 3385
rect 1374 3365 1544 3375
rect 1864 3365 2104 3375
rect 2464 3365 2974 3375
rect 1354 3355 1544 3365
rect 1894 3355 2104 3365
rect 2484 3355 2964 3365
rect 1324 3345 1544 3355
rect 1904 3345 2094 3355
rect 1314 3335 1544 3345
rect 1914 3335 2094 3345
rect 2504 3345 2954 3355
rect 2504 3335 2944 3345
rect 1284 3325 1544 3335
rect 1944 3325 2084 3335
rect 1264 3315 1544 3325
rect 1954 3315 2084 3325
rect 2514 3325 2924 3335
rect 2514 3315 2914 3325
rect 1254 3305 1554 3315
rect 1234 3295 1554 3305
rect 1954 3305 2074 3315
rect 1954 3295 2034 3305
rect 2524 3295 2904 3315
rect 1214 3285 1554 3295
rect 1964 3285 2024 3295
rect 2524 3285 2894 3295
rect 1194 3275 1564 3285
rect 1994 3275 2004 3285
rect 2514 3275 2884 3285
rect 1174 3265 1574 3275
rect 2504 3265 2874 3275
rect 1154 3255 1584 3265
rect 2494 3255 2864 3265
rect 1134 3245 1594 3255
rect 2484 3245 2854 3255
rect 1104 3235 1594 3245
rect 2364 3235 2374 3245
rect 2454 3235 2854 3245
rect 1084 3225 1604 3235
rect 2354 3225 2384 3235
rect 1064 3215 1614 3225
rect 2364 3215 2384 3225
rect 2434 3225 2844 3235
rect 1044 3205 1614 3215
rect 2434 3205 2834 3225
rect 1024 3195 1624 3205
rect 2434 3195 2824 3205
rect 994 3185 1634 3195
rect 2364 3185 2414 3195
rect 2424 3185 2824 3195
rect 974 3175 1644 3185
rect 2364 3175 2814 3185
rect 944 3165 1654 3175
rect 2364 3165 2804 3175
rect 904 3155 1654 3165
rect 2404 3155 2804 3165
rect 874 3145 1664 3155
rect 2404 3145 2794 3155
rect 3724 3145 3754 3155
rect 844 3135 1674 3145
rect 2394 3135 2784 3145
rect 3724 3135 3734 3145
rect 814 3125 1694 3135
rect 784 3115 1704 3125
rect 2394 3115 2774 3135
rect 744 3105 1714 3115
rect 2394 3105 2764 3115
rect 694 3095 1724 3105
rect 2404 3095 2754 3105
rect 654 3085 1744 3095
rect 604 3075 1754 3085
rect 2404 3075 2744 3095
rect 574 3065 1764 3075
rect 2404 3065 2734 3075
rect 544 3055 1774 3065
rect 515 3045 1774 3055
rect 2404 3055 2724 3065
rect 2404 3045 2714 3055
rect 515 3035 1784 3045
rect 2414 3035 2714 3045
rect 515 3025 1804 3035
rect 2424 3025 2714 3035
rect 515 3015 1814 3025
rect 515 3005 1834 3015
rect 2224 3005 2264 3015
rect 2434 3005 2464 3025
rect 2484 3005 2704 3025
rect 515 2995 1854 3005
rect 515 2985 1864 2995
rect 2214 2985 2274 3005
rect 2414 2995 2694 3005
rect 515 2975 1884 2985
rect 2204 2975 2274 2985
rect 2404 2985 2694 2995
rect 515 2965 1894 2975
rect 2214 2965 2264 2975
rect 515 2955 1904 2965
rect 2234 2955 2254 2965
rect 2404 2955 2684 2985
rect 515 2945 1924 2955
rect 2394 2945 2684 2955
rect 515 2935 1944 2945
rect 2384 2935 2684 2945
rect 515 2925 1954 2935
rect 2374 2925 2674 2935
rect 515 2915 1984 2925
rect 2364 2915 2674 2925
rect 515 2905 2014 2915
rect 2174 2905 2194 2915
rect 2354 2905 2674 2915
rect 515 2895 2024 2905
rect 515 2885 2034 2895
rect 2164 2885 2214 2905
rect 2344 2895 2684 2905
rect 2324 2885 2684 2895
rect 515 2875 2054 2885
rect 2104 2875 2214 2885
rect 2294 2875 2674 2885
rect 515 2835 2224 2875
rect 2274 2865 2674 2875
rect 2264 2855 2674 2865
rect 515 2815 2214 2835
rect 515 2805 2224 2815
rect 515 2795 2234 2805
rect 2264 2795 2684 2855
rect 515 2765 2684 2795
rect 515 2755 2294 2765
rect 2324 2755 2684 2765
rect 515 2745 2684 2755
rect 515 2675 2694 2745
rect 4044 2715 4094 2725
rect 4034 2705 4124 2715
rect 4024 2695 4134 2705
rect 4014 2685 4154 2695
rect 4004 2675 4164 2685
rect 515 2605 2684 2675
rect 3994 2665 4184 2675
rect 3974 2655 4194 2665
rect 3964 2645 4204 2655
rect 3944 2635 4224 2645
rect 3924 2625 4244 2635
rect 3914 2615 4254 2625
rect 3894 2605 4274 2615
rect 515 2565 2674 2605
rect 3884 2595 4294 2605
rect 3874 2585 4298 2595
rect 3864 2575 4298 2585
rect 3854 2565 4298 2575
rect 515 2495 2664 2565
rect 3844 2545 4298 2565
rect 3834 2535 4298 2545
rect 3824 2525 4298 2535
rect 3814 2515 4298 2525
rect 3804 2505 4298 2515
rect 515 2465 2654 2495
rect 3794 2475 4298 2505
rect 515 2425 2644 2465
rect 3784 2455 4298 2475
rect 3774 2435 4298 2455
rect 3734 2425 3744 2435
rect 3764 2425 4298 2435
rect 515 2385 2634 2425
rect 3724 2415 4298 2425
rect 3714 2405 4298 2415
rect 515 2355 2624 2385
rect 3704 2375 4298 2405
rect 3694 2355 4298 2375
rect 515 2315 2614 2355
rect 3684 2345 4298 2355
rect 3674 2325 4298 2345
rect 515 2285 2604 2315
rect 3664 2305 4298 2325
rect 3654 2295 4298 2305
rect 3644 2285 4298 2295
rect 515 2265 2594 2285
rect 3634 2275 4298 2285
rect 3624 2265 4298 2275
rect 515 2235 2584 2265
rect 3614 2245 4298 2265
rect 3604 2235 4298 2245
rect 515 2215 2574 2235
rect 3594 2215 4298 2235
rect 515 2205 2564 2215
rect 515 2185 2554 2205
rect 3584 2195 4298 2215
rect 3574 2185 4298 2195
rect 515 2175 2544 2185
rect 3564 2175 4298 2185
rect 515 2155 2534 2175
rect 3554 2165 4298 2175
rect 3544 2155 4298 2165
rect 515 2135 2524 2155
rect 3534 2145 4298 2155
rect 3524 2135 4298 2145
rect 515 2115 2514 2135
rect 3514 2125 4298 2135
rect 3504 2115 4298 2125
rect 515 2095 2504 2115
rect 3494 2095 4298 2115
rect 515 2085 2494 2095
rect 3474 2085 4298 2095
rect 515 2065 2484 2085
rect 3464 2075 4298 2085
rect 3454 2065 4298 2075
rect 515 2055 2474 2065
rect 3434 2055 4298 2065
rect 515 2025 2464 2055
rect 3424 2045 4298 2055
rect 3404 2035 4298 2045
rect 515 2005 2454 2025
rect 3394 2015 4298 2035
rect 3384 2005 4298 2015
rect 515 1985 2444 2005
rect 3374 1995 4298 2005
rect 3364 1985 4298 1995
rect 515 1965 2434 1985
rect 3354 1975 4298 1985
rect 3344 1965 4298 1975
rect 515 1955 2424 1965
rect 3334 1955 4298 1965
rect 515 1935 2414 1955
rect 3324 1945 4298 1955
rect 3314 1935 4298 1945
rect 515 1915 2404 1935
rect 515 1905 2394 1915
rect 3304 1905 4298 1935
rect 515 1885 2384 1905
rect 3294 1885 4298 1905
rect 515 1875 2374 1885
rect 515 1855 2364 1875
rect 3284 1865 4298 1885
rect 515 1845 2354 1855
rect 3274 1845 4298 1865
rect 515 1825 2344 1845
rect 3264 1835 4298 1845
rect 515 1805 2334 1825
rect 3254 1815 4298 1835
rect 3244 1805 4298 1815
rect 515 1785 2324 1805
rect 3234 1795 4298 1805
rect 3224 1785 4298 1795
rect 515 1765 2314 1785
rect 3214 1775 4298 1785
rect 3204 1765 4298 1775
rect 515 1745 2304 1765
rect 3194 1745 4298 1765
rect 515 1725 2294 1745
rect 3184 1735 4298 1745
rect 515 1705 2284 1725
rect 3174 1715 4298 1735
rect 3164 1705 4298 1715
rect 515 1685 2274 1705
rect 3154 1685 4298 1705
rect 515 1665 2264 1685
rect 3144 1665 4298 1685
rect 515 1645 2254 1665
rect 3134 1655 4298 1665
rect 515 1625 2244 1645
rect 515 1605 2234 1625
rect 3124 1615 4298 1655
rect 3114 1605 3254 1615
rect 3304 1605 4298 1615
rect 515 1585 2224 1605
rect 3114 1595 3244 1605
rect 3314 1595 4298 1605
rect 3104 1585 3234 1595
rect 3324 1585 4298 1595
rect 515 1565 2214 1585
rect 3104 1575 3224 1585
rect 3344 1575 4298 1585
rect 3094 1565 3214 1575
rect 3354 1565 4298 1575
rect 515 1545 2204 1565
rect 3094 1555 3204 1565
rect 3364 1555 4298 1565
rect 3094 1545 3194 1555
rect 3384 1545 4298 1555
rect 515 1525 2194 1545
rect 3094 1535 3184 1545
rect 3394 1535 4298 1545
rect 3084 1525 3174 1535
rect 3404 1525 4298 1535
rect 515 1505 2184 1525
rect 3084 1515 3164 1525
rect 3414 1515 4298 1525
rect 3074 1505 3154 1515
rect 3424 1505 4298 1515
rect 515 1485 2174 1505
rect 3074 1495 3144 1505
rect 3434 1495 4298 1505
rect 3074 1485 3134 1495
rect 3444 1485 4298 1495
rect 515 1465 2164 1485
rect 3064 1475 3114 1485
rect 3454 1475 4298 1485
rect 3064 1465 3104 1475
rect 3464 1465 4298 1475
rect 515 1445 2154 1465
rect 3064 1455 3084 1465
rect 3474 1455 4298 1465
rect 3484 1445 4298 1455
rect 515 1425 2144 1445
rect 3494 1425 4298 1445
rect 515 1395 2134 1425
rect 3504 1415 4298 1425
rect 3514 1405 4298 1415
rect 3534 1395 4298 1405
rect 515 1375 2124 1395
rect 3544 1385 4298 1395
rect 3554 1375 4298 1385
rect 515 1355 2114 1375
rect 3564 1365 4298 1375
rect 3574 1355 4298 1365
rect 515 1335 2104 1355
rect 3584 1345 4298 1355
rect 515 1315 2094 1335
rect 3594 1325 4298 1345
rect 3604 1315 4298 1325
rect 515 1305 2084 1315
rect 3614 1305 4298 1315
rect 515 1285 2074 1305
rect 3624 1295 4298 1305
rect 515 1275 2064 1285
rect 3634 1275 4298 1295
rect 515 1255 2054 1275
rect 3644 1265 4298 1275
rect 515 1235 2044 1255
rect 3654 1245 4298 1265
rect 515 1215 2034 1235
rect 3664 1225 4298 1245
rect 2974 1215 3024 1225
rect 515 1195 2024 1215
rect 2964 1205 3054 1215
rect 3674 1205 4298 1225
rect 2954 1195 3064 1205
rect 515 1185 2014 1195
rect 2954 1185 3084 1195
rect 515 1165 2004 1185
rect 2944 1175 3094 1185
rect 2944 1165 3104 1175
rect 515 1145 1994 1165
rect 2934 1155 3124 1165
rect 3684 1155 4298 1205
rect 2934 1145 3144 1155
rect 515 1135 1984 1145
rect 2934 1135 3154 1145
rect 3674 1135 4298 1155
rect 515 1115 1974 1135
rect 2934 1125 3164 1135
rect 2934 1115 3184 1125
rect 3664 1115 4298 1135
rect 515 1095 1964 1115
rect 2924 1105 3194 1115
rect 3654 1105 4298 1115
rect 2924 1095 3214 1105
rect 3644 1095 4298 1105
rect 515 1085 1954 1095
rect 2924 1085 3224 1095
rect 515 1065 1944 1085
rect 2914 1075 3244 1085
rect 3634 1075 4298 1095
rect 2914 1065 3264 1075
rect 3624 1065 4298 1075
rect 515 1045 1934 1065
rect 2904 1055 3284 1065
rect 2904 1045 3294 1055
rect 3614 1045 4298 1065
rect 515 1035 1924 1045
rect 2894 1035 3314 1045
rect 3604 1035 4298 1045
rect 515 1015 1914 1035
rect 2894 1025 3334 1035
rect 3594 1025 4298 1035
rect 2884 1015 3344 1025
rect 3584 1015 4298 1025
rect 515 995 1904 1015
rect 2884 1005 3354 1015
rect 3574 1005 4298 1015
rect 2884 995 3374 1005
rect 3564 995 4298 1005
rect 515 985 1894 995
rect 2874 985 3384 995
rect 3554 985 4298 995
rect 515 965 1884 985
rect 2874 975 3394 985
rect 3544 975 4298 985
rect 2874 965 3404 975
rect 3534 965 4298 975
rect 515 955 1874 965
rect 2874 955 3424 965
rect 3514 955 4298 965
rect 515 935 1864 955
rect 2864 945 3444 955
rect 3504 945 4298 955
rect 2864 935 3454 945
rect 3494 935 4298 945
rect 515 925 1854 935
rect 515 905 1844 925
rect 2854 915 3454 935
rect 3474 925 4298 935
rect 3464 915 4298 925
rect 2854 905 3444 915
rect 515 895 1834 905
rect 2844 895 3434 905
rect 3474 895 4298 915
rect 515 875 1824 895
rect 2844 885 3414 895
rect 3484 885 4298 895
rect 2844 875 3404 885
rect 3504 875 4298 885
rect 515 865 1814 875
rect 2834 865 3384 875
rect 3524 865 4298 875
rect 515 855 1804 865
rect 2834 855 3374 865
rect 3534 855 4298 865
rect 515 835 1794 855
rect 2834 845 3364 855
rect 3544 845 4298 855
rect 2824 835 3344 845
rect 3554 835 4298 845
rect 515 815 1784 835
rect 2824 825 3334 835
rect 3564 825 4298 835
rect 2814 815 3324 825
rect 3574 815 4298 825
rect 515 805 1774 815
rect 2814 805 3304 815
rect 3584 805 4298 815
rect 515 785 1764 805
rect 2814 795 3294 805
rect 3604 795 4298 805
rect 2804 785 3274 795
rect 3614 785 4298 795
rect 515 775 1754 785
rect 2804 775 3264 785
rect 3624 775 4298 785
rect 515 765 1744 775
rect 2794 765 3254 775
rect 515 755 1734 765
rect 2794 755 3234 765
rect 3634 755 4298 775
rect 515 735 1724 755
rect 2794 745 3224 755
rect 3644 745 4298 755
rect 2784 735 3214 745
rect 3654 735 4298 745
rect 515 715 1714 735
rect 2774 725 3194 735
rect 3664 725 4298 735
rect 2774 715 3174 725
rect 3674 715 4298 725
rect 515 705 1704 715
rect 2774 705 3164 715
rect 3684 705 4298 715
rect 515 695 1694 705
rect 2774 695 2794 705
rect 2834 695 3144 705
rect 3694 695 4298 705
rect 515 675 1684 695
rect 2844 685 3134 695
rect 3704 685 4298 695
rect 2864 675 3114 685
rect 3714 675 4298 685
rect 515 665 1674 675
rect 2874 665 3104 675
rect 3724 665 4298 675
rect 515 655 1664 665
rect 2884 655 3084 665
rect 515 645 1654 655
rect 2894 645 3074 655
rect 3734 645 4298 665
rect 515 625 1644 645
rect 2904 635 3054 645
rect 2914 625 3044 635
rect 515 615 1634 625
rect 2914 615 3034 625
rect 515 595 1624 615
rect 2924 605 3024 615
rect 2934 595 3014 605
rect 515 585 1614 595
rect 2944 585 2994 595
rect 515 575 1604 585
rect 2954 575 2984 585
rect 515 565 1594 575
rect 515 555 1584 565
rect 515 545 754 555
rect 1034 545 1574 555
rect 515 535 644 545
rect 1094 535 1564 545
rect 3744 535 4298 645
rect 515 525 584 535
rect 1144 525 1554 535
rect 3734 525 4298 535
rect 515 515 544 525
rect 1174 515 1544 525
rect 1204 505 1534 515
rect 3724 505 4298 525
rect 1234 495 1524 505
rect 2964 495 2984 505
rect 3714 495 4298 505
rect 1254 485 1524 495
rect 1274 475 1514 485
rect 2944 475 2994 495
rect 3704 485 4298 495
rect 3694 475 4298 485
rect 1284 465 1494 475
rect 2934 465 2994 475
rect 3684 465 4298 475
rect 1294 455 1484 465
rect 2924 455 2994 465
rect 3674 455 4298 465
rect 1304 435 1474 455
rect 2914 445 2984 455
rect 3664 445 4298 455
rect 2914 435 2974 445
rect 3654 435 4298 445
rect 1314 425 1464 435
rect 2904 425 2974 435
rect 3634 425 4298 435
rect 1324 415 1454 425
rect 2904 415 2954 425
rect 3014 415 3024 425
rect 3624 415 4298 425
rect 1324 405 1444 415
rect 2894 405 2944 415
rect 3004 405 3034 415
rect 3614 405 4298 415
rect 1324 395 1434 405
rect 2884 395 2944 405
rect 3014 395 3044 405
rect 3594 395 4298 405
rect 1334 385 1424 395
rect 1334 375 1414 385
rect 2874 375 2934 395
rect 3014 385 3054 395
rect 3584 385 4298 395
rect 3024 375 3054 385
rect 3574 375 4298 385
rect 1334 365 1394 375
rect 2864 365 2924 375
rect 3564 365 4298 375
rect 1354 355 1364 365
rect 2854 355 2914 365
rect 3554 355 4298 365
rect 2844 345 2904 355
rect 3544 345 4298 355
rect 2834 335 2894 345
rect 3524 335 4298 345
rect 2824 325 2884 335
rect 3514 325 4298 335
rect 2814 315 2884 325
rect 3494 315 4298 325
rect 2804 305 2864 315
rect 3484 305 4298 315
rect 2794 295 2864 305
rect 3134 295 3144 305
rect 3474 295 4298 305
rect 2794 285 2854 295
rect 3134 285 3154 295
rect 3454 285 4298 295
rect 2784 275 2844 285
rect 3144 275 3154 285
rect 3434 275 4298 285
rect 2774 265 2834 275
rect 3424 265 4298 275
rect 2764 255 2824 265
rect 3404 255 4298 265
rect 2754 245 2814 255
rect 3174 245 3194 255
rect 3394 245 4298 255
rect 2744 235 2804 245
rect 3184 235 3204 245
rect 3374 235 4298 245
rect 2734 225 2794 235
rect 3194 225 3214 235
rect 3354 225 4298 235
rect 2724 215 2784 225
rect 3204 215 3234 225
rect 3344 215 4298 225
rect 2714 205 2774 215
rect 3214 205 3254 215
rect 3324 205 4298 215
rect 2574 195 2644 205
rect 2704 195 2764 205
rect 3224 195 3274 205
rect 3294 195 3424 205
rect 2574 185 2664 195
rect 2694 185 2754 195
rect 3234 185 3404 195
rect 2564 175 2744 185
rect 3244 175 3394 185
rect 3464 175 4298 205
rect 2574 165 2734 175
rect 3254 165 3374 175
rect 2604 155 2724 165
rect 3254 155 3354 165
rect 2624 145 2724 155
rect 3264 145 3344 155
rect 3454 145 4298 175
rect 2634 135 2714 145
rect 3274 135 3324 145
rect 2644 125 2704 135
rect 3284 125 3304 135
rect 2654 115 2684 125
rect 3444 115 4298 145
rect 3434 95 4298 115
rect 3414 85 4298 95
rect 3404 75 4298 85
rect 3394 65 4298 75
rect 3374 55 4298 65
rect 3364 45 4298 55
rect 2514 35 2564 45
rect 3354 35 4298 45
rect 2504 25 2584 35
rect 3334 25 4298 35
rect 2494 15 2604 25
rect 3324 15 4298 25
rect 2494 5 2614 15
rect 3314 5 4298 15
rect 2484 -5 2634 5
rect 3304 -3 4298 5
rect 3304 -5 4514 -3
rect 2484 -15 2654 -5
rect 3294 -15 4514 -5
use erin-threshold  erin-threshold_0
timestamp 1419146600
transform 1 0 3197 0 1 -721
box 1134 718 4724 7241
<< end >>
