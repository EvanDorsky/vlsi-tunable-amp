magic
tech scmos
timestamp 1421379733
<< nwell >>
rect 766 603 770 607
rect 766 599 769 600
rect 766 579 770 583
rect 518 511 562 514
rect 636 511 670 514
rect 162 258 196 511
<< pwell >>
rect -7 511 481 663
rect 553 648 585 668
rect 1285 663 1589 667
rect 753 618 756 619
rect 761 613 762 614
rect 759 612 762 613
rect 759 611 761 612
rect 760 608 761 611
rect 752 604 753 607
rect 760 597 763 608
rect 953 514 1589 663
rect -7 258 162 511
rect -7 255 179 258
rect -7 247 178 255
rect -7 242 170 247
<< electrodecontact >>
rect 151 437 155 629
rect 468 522 472 636
rect 982 525 986 643
rect 1298 525 1302 643
rect 1686 268 1690 420
<< electrodecap >>
rect 1 435 157 631
rect 194 520 474 642
rect 980 523 1259 649
rect 1296 523 1575 649
<< psubstratepcontact >>
rect -4 639 162 643
rect 182 515 186 647
rect 1267 518 1271 654
rect 1284 518 1288 654
<< polysilicon >>
rect -4 430 162 633
rect 192 515 479 647
rect 975 518 1261 654
rect 1294 518 1580 654
<< polycontact >>
rect -4 633 162 637
rect 188 515 192 647
rect 865 518 869 522
rect 1261 518 1265 654
rect 1290 518 1294 654
<< metal1 >>
rect 883 691 885 692
rect 865 688 885 691
rect 167 680 266 684
rect -4 637 162 639
rect 167 589 171 680
rect 266 654 269 669
rect 865 668 869 688
rect 838 661 862 664
rect 1238 661 1242 669
rect 762 659 1242 661
rect 762 657 844 659
rect 858 657 1242 659
rect 545 654 593 655
rect 266 652 775 654
rect 266 651 548 652
rect 590 651 771 652
rect 155 585 171 589
rect 186 515 188 647
rect 753 618 756 619
rect 735 520 790 524
rect 1265 518 1267 654
rect 1288 518 1290 654
rect 1686 420 1689 674
<< m2contact >>
rect 889 673 893 677
rect 473 664 477 668
rect 480 664 484 668
rect 865 664 869 668
rect 1238 669 1242 673
rect 758 657 762 661
rect 771 648 775 652
rect 982 643 986 647
rect 468 636 472 640
rect 823 625 827 629
rect 766 603 770 607
rect 766 579 770 583
rect 766 555 770 559
rect 766 531 770 535
rect 865 522 869 526
rect 1298 643 1302 647
<< metal2 >>
rect 765 673 889 674
rect 893 673 986 677
rect 765 671 892 673
rect 468 664 473 668
rect 561 667 577 668
rect 484 665 749 667
rect 484 664 564 665
rect 574 664 749 665
rect 468 640 472 664
rect 746 636 749 664
rect 746 633 756 636
rect 753 607 756 633
rect 759 614 762 657
rect 765 620 768 671
rect 771 626 774 648
rect 777 629 786 633
rect 771 623 776 626
rect 782 625 823 629
rect 765 617 770 620
rect 759 611 763 614
rect 752 604 756 607
rect 752 576 755 604
rect 760 600 763 611
rect 767 607 770 617
rect 760 597 769 600
rect 766 583 769 597
rect 752 573 769 576
rect 766 559 769 573
rect 773 535 776 623
rect 770 532 776 535
rect 865 526 869 664
rect 982 647 986 673
rect 1242 669 1302 673
rect 1298 647 1302 669
use resistors  resistors_0
timestamp 1419289491
transform -1 0 1688 0 -1 699
box -21 -26 1675 36
use spi-interface  spi-interface_0
timestamp 1419262457
transform 0 1 502 -1 0 622
box -27 -21 108 279
use amplifier  amplifier_0
timestamp 1419285127
transform 1 0 0 0 1 0
box 0 0 1733 655
<< labels >>
rlabel metal2 765 634 768 636 1 B0
rlabel metal2 759 634 762 636 1 B1
rlabel metal2 753 634 756 636 1 B2
rlabel metal2 771 634 774 636 1 B3
<< end >>
