magic
tech scmos
magscale 1 3
timestamp 1419061922
<< metal1 >>
rect 3220 7190 3250 7200
rect 3180 7180 3280 7190
rect 3140 7170 3300 7180
rect 3120 7160 3320 7170
rect 3100 7150 3330 7160
rect 3080 7140 3340 7150
rect 3070 7130 3450 7140
rect 3070 7120 3460 7130
rect 3080 7110 3480 7120
rect 3080 7100 3490 7110
rect 2950 7090 2970 7100
rect 3080 7090 3510 7100
rect 2940 7080 2990 7090
rect 3080 7080 3540 7090
rect 2790 7070 2820 7080
rect 2780 7060 2820 7070
rect 2940 7060 3010 7080
rect 3080 7070 3560 7080
rect 3070 7060 3570 7070
rect 2770 7050 2810 7060
rect 2750 7040 2810 7050
rect 2950 7050 3010 7060
rect 3060 7050 3580 7060
rect 3690 7050 3720 7060
rect 2950 7040 3020 7050
rect 3050 7040 3610 7050
rect 3670 7040 3760 7050
rect 3820 7040 3890 7050
rect 2740 7030 2810 7040
rect 2960 7030 3900 7040
rect 2720 7020 2860 7030
rect 2960 7020 3910 7030
rect 2700 7010 2860 7020
rect 2670 7000 2860 7010
rect 2650 6990 2860 7000
rect 2640 6980 2860 6990
rect 2990 7010 3950 7020
rect 4050 7010 4160 7020
rect 2990 7000 3960 7010
rect 4030 7000 4170 7010
rect 2990 6990 3980 7000
rect 3990 6990 4160 7000
rect 2990 6980 4160 6990
rect 2650 6960 2850 6980
rect 2970 6970 4150 6980
rect 2950 6960 4150 6970
rect 4410 6960 4450 6970
rect 2590 6950 2600 6960
rect 2580 6940 2600 6950
rect 2570 6920 2600 6940
rect 2660 6950 2850 6960
rect 2940 6950 4150 6960
rect 4400 6950 4460 6960
rect 2660 6940 2890 6950
rect 2920 6940 4150 6950
rect 2660 6930 4150 6940
rect 2660 6920 4160 6930
rect 4250 6920 4260 6930
rect 2560 6900 2590 6920
rect 2650 6910 2810 6920
rect 2820 6910 4370 6920
rect 2640 6900 2780 6910
rect 2840 6900 4380 6910
rect 2550 6890 2590 6900
rect 2630 6890 2780 6900
rect 2560 6880 2590 6890
rect 2620 6880 2790 6890
rect 2850 6880 4390 6900
rect 2550 6870 2800 6880
rect 2840 6870 4100 6880
rect 4110 6870 4400 6880
rect 2520 6860 4090 6870
rect 2490 6850 4090 6860
rect 4110 6850 4410 6870
rect 2450 6840 4020 6850
rect 4110 6840 4420 6850
rect 2450 6830 4000 6840
rect 4100 6830 4420 6840
rect 2440 6820 4000 6830
rect 4090 6820 4420 6830
rect 2430 6810 4020 6820
rect 4080 6810 4430 6820
rect 4610 6810 4660 6820
rect 2430 6800 3680 6810
rect 3720 6800 4430 6810
rect 4570 6800 4670 6810
rect 2420 6790 3670 6800
rect 2410 6780 3660 6790
rect 3720 6780 4440 6800
rect 4550 6790 4680 6800
rect 4550 6780 4690 6790
rect 2350 6770 3260 6780
rect 3270 6770 3480 6780
rect 3490 6770 3650 6780
rect 2330 6750 3250 6770
rect 3270 6760 3460 6770
rect 3500 6760 3650 6770
rect 3720 6760 4450 6780
rect 4540 6770 4710 6780
rect 4540 6760 4720 6770
rect 3270 6750 3450 6760
rect 3490 6750 3650 6760
rect 3710 6750 4470 6760
rect 4540 6750 4730 6760
rect 2320 6740 3250 6750
rect 3280 6740 3450 6750
rect 3480 6740 4480 6750
rect 4540 6740 4740 6750
rect 2320 6730 3260 6740
rect 3270 6730 3440 6740
rect 3470 6730 4490 6740
rect 4540 6730 4750 6740
rect 2320 6720 3300 6730
rect 3340 6720 3440 6730
rect 3460 6720 4500 6730
rect 4540 6720 4760 6730
rect 2320 6710 3290 6720
rect 3340 6710 3430 6720
rect 3450 6710 4510 6720
rect 4530 6710 4760 6720
rect 2320 6690 3280 6710
rect 3340 6700 3420 6710
rect 3330 6690 3420 6700
rect 3450 6700 3660 6710
rect 3690 6700 4770 6710
rect 2310 6680 3270 6690
rect 3320 6680 3410 6690
rect 2310 6670 3250 6680
rect 3320 6670 3390 6680
rect 3450 6670 3650 6700
rect 3700 6680 4780 6700
rect 3700 6670 4790 6680
rect 2290 6660 3230 6670
rect 3320 6660 3370 6670
rect 2280 6650 3220 6660
rect 2270 6640 3140 6650
rect 3190 6640 3210 6650
rect 3320 6640 3360 6660
rect 3440 6650 3650 6670
rect 3690 6660 4780 6670
rect 3690 6650 4400 6660
rect 4430 6650 4790 6660
rect 4820 6650 4830 6660
rect 3430 6640 3660 6650
rect 3680 6640 4400 6650
rect 4450 6640 4840 6650
rect 2250 6630 3100 6640
rect 3310 6630 3360 6640
rect 3420 6630 4390 6640
rect 2250 6620 3080 6630
rect 3300 6620 3370 6630
rect 3410 6620 3930 6630
rect 3960 6620 4390 6630
rect 4460 6630 4840 6640
rect 4460 6620 4680 6630
rect 4710 6620 4840 6630
rect 2240 6610 3070 6620
rect 3200 6610 3210 6620
rect 3290 6610 3920 6620
rect 3960 6610 4400 6620
rect 4440 6610 4670 6620
rect 4720 6610 4830 6620
rect 2230 6600 3070 6610
rect 3190 6600 3220 6610
rect 3280 6600 3910 6610
rect 3950 6600 4400 6610
rect 4420 6600 4600 6610
rect 2220 6590 3080 6600
rect 3180 6590 3230 6600
rect 3260 6590 3900 6600
rect 3940 6590 4600 6600
rect 4610 6600 4650 6610
rect 4760 6600 4810 6610
rect 4610 6590 4640 6600
rect 2220 6580 3130 6590
rect 3170 6580 3890 6590
rect 3920 6580 4640 6590
rect 2220 6570 3880 6580
rect 3900 6570 4630 6580
rect 2220 6550 3620 6570
rect 3640 6560 3870 6570
rect 3890 6560 4640 6570
rect 3650 6550 4640 6560
rect 2220 6540 3610 6550
rect 2230 6520 3610 6540
rect 3650 6530 4650 6550
rect 3640 6520 4650 6530
rect 4800 6540 4830 6550
rect 4800 6520 4840 6540
rect 2230 6510 2670 6520
rect 2700 6510 4660 6520
rect 4800 6510 4850 6520
rect 2230 6500 2660 6510
rect 2710 6500 3060 6510
rect 3080 6500 4660 6510
rect 4790 6500 4850 6510
rect 2230 6490 2590 6500
rect 2640 6490 2650 6500
rect 2710 6490 3050 6500
rect 3080 6490 4670 6500
rect 2230 6480 2580 6490
rect 2230 6450 2570 6480
rect 2610 6460 2650 6470
rect 2720 6460 3040 6490
rect 3080 6480 3480 6490
rect 3490 6480 4680 6490
rect 4780 6480 4850 6500
rect 3070 6460 3480 6480
rect 3500 6460 4700 6480
rect 4790 6460 4850 6480
rect 2580 6450 2660 6460
rect 2240 6440 2660 6450
rect 2730 6450 3050 6460
rect 3060 6450 3780 6460
rect 2730 6440 3780 6450
rect 3810 6440 4710 6460
rect 4780 6440 4850 6460
rect 2250 6420 2670 6440
rect 2730 6430 2980 6440
rect 3020 6430 3780 6440
rect 3800 6430 4710 6440
rect 4760 6430 4850 6440
rect 2250 6410 2530 6420
rect 2570 6410 2670 6420
rect 2720 6410 2980 6430
rect 3010 6420 4710 6430
rect 4750 6420 4850 6430
rect 3000 6410 4830 6420
rect 2250 6400 2510 6410
rect 2580 6400 2670 6410
rect 2240 6390 2500 6400
rect 2570 6390 2680 6400
rect 2710 6390 4820 6410
rect 4830 6390 4860 6400
rect 4950 6390 5010 6400
rect 2240 6380 2490 6390
rect 2560 6380 4870 6390
rect 4940 6380 5020 6390
rect 2240 6370 2480 6380
rect 2550 6370 4890 6380
rect 4930 6370 5020 6380
rect 2230 6360 2720 6370
rect 2760 6360 5020 6370
rect 2230 6350 2700 6360
rect 2220 6340 2590 6350
rect 2640 6340 2690 6350
rect 2770 6340 5020 6360
rect 2210 6330 2580 6340
rect 2200 6320 2570 6330
rect 2760 6320 5020 6340
rect 2130 6310 2150 6320
rect 2190 6310 2560 6320
rect 2750 6310 5020 6320
rect 2100 6300 2550 6310
rect 2090 6290 2540 6300
rect 2750 6290 5010 6310
rect 2080 6280 2530 6290
rect 2740 6280 5010 6290
rect 2070 6270 2530 6280
rect 2630 6270 2650 6280
rect 2720 6270 3630 6280
rect 3670 6270 3800 6280
rect 3850 6270 5020 6280
rect 2050 6260 2540 6270
rect 2550 6260 2660 6270
rect 2710 6260 3620 6270
rect 3680 6260 3770 6270
rect 2040 6250 3620 6260
rect 3690 6250 3770 6260
rect 2020 6240 3620 6250
rect 2010 6230 3620 6240
rect 3700 6230 3770 6250
rect 3860 6260 5030 6270
rect 3860 6250 4850 6260
rect 4860 6250 5030 6260
rect 3860 6240 4830 6250
rect 4870 6240 5040 6250
rect 3850 6230 4830 6240
rect 2000 6220 3630 6230
rect 3700 6220 3750 6230
rect 3830 6220 4830 6230
rect 4880 6220 5040 6240
rect 1910 6210 1940 6220
rect 2000 6210 3740 6220
rect 3820 6210 4830 6220
rect 1900 6200 1950 6210
rect 1890 6190 1950 6200
rect 2000 6200 3730 6210
rect 1890 6180 1940 6190
rect 1880 6160 1940 6180
rect 2000 6180 3740 6200
rect 3810 6190 4830 6210
rect 3810 6180 4410 6190
rect 4420 6180 4840 6190
rect 2000 6170 3750 6180
rect 3810 6170 4840 6180
rect 1990 6160 3760 6170
rect 3800 6160 4840 6170
rect 4870 6160 5040 6220
rect 1880 6150 1920 6160
rect 1980 6150 4840 6160
rect 1880 6140 1910 6150
rect 1970 6130 4850 6150
rect 4880 6140 5040 6160
rect 1960 6120 3550 6130
rect 3560 6120 4850 6130
rect 1960 6110 3520 6120
rect 3580 6110 4850 6120
rect 1960 6100 3500 6110
rect 3590 6100 4850 6110
rect 1950 6090 3490 6100
rect 3600 6090 4850 6100
rect 1950 6070 3480 6090
rect 1950 6060 3470 6070
rect 1950 6040 3480 6060
rect 1940 6030 3480 6040
rect 3590 6050 4850 6090
rect 4890 6110 5040 6140
rect 4890 6090 5030 6110
rect 4890 6080 5020 6090
rect 4900 6070 4960 6080
rect 4910 6060 4950 6070
rect 4930 6050 4940 6060
rect 3590 6040 4000 6050
rect 4040 6040 4840 6050
rect 3590 6030 3990 6040
rect 4080 6030 4840 6040
rect 1930 6020 3480 6030
rect 1870 6010 3480 6020
rect 3600 6010 3980 6030
rect 4110 6020 4840 6030
rect 4130 6010 4830 6020
rect 1860 5990 3490 6010
rect 3600 6000 3970 6010
rect 4140 6000 4830 6010
rect 1860 5980 3500 5990
rect 3610 5980 3970 6000
rect 4120 5990 4930 6000
rect 4080 5980 5000 5990
rect 1850 5970 3500 5980
rect 1850 5960 3490 5970
rect 3600 5960 3960 5980
rect 4030 5970 5050 5980
rect 5140 5970 5170 5980
rect 4000 5960 5170 5970
rect 1850 5950 3480 5960
rect 3650 5950 3960 5960
rect 3970 5950 5170 5960
rect 1850 5940 3470 5950
rect 3660 5940 5160 5950
rect 1850 5930 3460 5940
rect 3670 5930 5160 5940
rect 1850 5920 3450 5930
rect 3680 5920 5150 5930
rect 1840 5900 3440 5920
rect 3700 5910 3740 5920
rect 3820 5910 5140 5920
rect 3840 5900 5130 5910
rect 1840 5890 3430 5900
rect 3820 5890 5110 5900
rect 1830 5880 3420 5890
rect 3800 5880 5080 5890
rect 1830 5870 3410 5880
rect 3780 5870 5030 5880
rect 1840 5860 3360 5870
rect 3760 5860 5010 5870
rect 1840 5850 3330 5860
rect 3740 5850 5000 5860
rect 1850 5840 3280 5850
rect 3720 5840 4990 5850
rect 1850 5830 3260 5840
rect 3710 5830 4980 5840
rect 1850 5820 3250 5830
rect 3690 5820 4980 5830
rect 1850 5810 3230 5820
rect 3680 5810 3910 5820
rect 3940 5810 4970 5820
rect 1840 5800 3210 5810
rect 3660 5800 3900 5810
rect 3950 5800 4970 5810
rect 1840 5780 3190 5800
rect 3650 5790 3890 5800
rect 3970 5790 4960 5800
rect 3670 5780 3870 5790
rect 3980 5780 4810 5790
rect 4850 5780 4960 5790
rect 1840 5770 3180 5780
rect 3680 5770 3810 5780
rect 3990 5770 4790 5780
rect 4880 5770 4960 5780
rect 1840 5760 3170 5770
rect 3690 5760 3760 5770
rect 4100 5760 4390 5770
rect 4450 5760 4760 5770
rect 4900 5760 4960 5770
rect 1830 5730 3170 5760
rect 3700 5750 3740 5760
rect 4110 5750 4380 5760
rect 4470 5750 4670 5760
rect 4120 5740 4360 5750
rect 4490 5740 4640 5750
rect 4130 5730 4340 5740
rect 4510 5730 4610 5740
rect 4910 5730 4960 5760
rect 1820 5720 3170 5730
rect 1810 5710 1920 5720
rect 1970 5710 3170 5720
rect 4150 5720 4320 5730
rect 4530 5720 4590 5730
rect 4150 5710 4270 5720
rect 4920 5710 4970 5730
rect 1800 5700 1860 5710
rect 1880 5700 1890 5710
rect 1800 5690 1820 5700
rect 2040 5690 3170 5710
rect 4160 5700 4250 5710
rect 4920 5700 4980 5710
rect 3530 5690 3570 5700
rect 4170 5690 4230 5700
rect 4930 5690 4980 5700
rect 1800 5680 1810 5690
rect 2040 5680 3180 5690
rect 3520 5680 3570 5690
rect 2040 5670 3190 5680
rect 3520 5670 3580 5680
rect 4930 5670 4990 5690
rect 2040 5660 3200 5670
rect 2030 5650 3210 5660
rect 3520 5650 3570 5670
rect 4940 5660 4990 5670
rect 2030 5640 3220 5650
rect 3520 5640 3560 5650
rect 4940 5640 4980 5660
rect 2020 5630 3230 5640
rect 2010 5620 3240 5630
rect 2000 5610 3240 5620
rect 2000 5600 3250 5610
rect 1990 5590 3250 5600
rect 1990 5580 3260 5590
rect 1980 5570 3260 5580
rect 3410 5570 3430 5580
rect 1970 5550 3270 5570
rect 3400 5560 3430 5570
rect 3390 5550 3430 5560
rect 1960 5540 3110 5550
rect 3130 5540 3280 5550
rect 3380 5540 3430 5550
rect 1960 5520 3100 5540
rect 3140 5530 3280 5540
rect 3370 5530 3420 5540
rect 3130 5520 3280 5530
rect 3360 5520 3420 5530
rect 1950 5500 3290 5520
rect 3350 5510 3420 5520
rect 3340 5500 3420 5510
rect 1950 5490 3320 5500
rect 3330 5490 3420 5500
rect 1940 5470 3430 5490
rect 1930 5460 3300 5470
rect 3310 5460 3440 5470
rect 1920 5440 3440 5460
rect 5240 5450 5290 5460
rect 5190 5440 5320 5450
rect 1910 5420 3440 5440
rect 4950 5430 5020 5440
rect 5150 5430 5330 5440
rect 4930 5420 5330 5430
rect 1900 5390 3440 5420
rect 4910 5410 5330 5420
rect 4900 5400 5330 5410
rect 4880 5390 5330 5400
rect 1900 5370 3450 5390
rect 4860 5380 5330 5390
rect 4850 5370 5330 5380
rect 1900 5360 3460 5370
rect 4830 5360 5330 5370
rect 1910 5350 3470 5360
rect 4810 5350 5330 5360
rect 1910 5340 3480 5350
rect 4800 5340 5330 5350
rect 1920 5330 3490 5340
rect 4780 5330 5330 5340
rect 1920 5320 3500 5330
rect 4760 5320 5320 5330
rect 1950 5310 3510 5320
rect 4740 5310 5320 5320
rect 1960 5300 3510 5310
rect 4720 5300 5190 5310
rect 5210 5300 5310 5310
rect 1970 5290 3520 5300
rect 4700 5290 5180 5300
rect 5220 5290 5310 5300
rect 1980 5270 3520 5290
rect 4300 5280 4410 5290
rect 4460 5280 4500 5290
rect 4680 5280 5180 5290
rect 4280 5270 4560 5280
rect 4660 5270 5180 5280
rect 1990 5260 3520 5270
rect 4240 5260 4610 5270
rect 4640 5260 5180 5270
rect 1990 5240 3510 5260
rect 4220 5250 5180 5260
rect 4200 5240 5180 5250
rect 5230 5240 5300 5290
rect 1990 5210 3500 5240
rect 4160 5230 5170 5240
rect 4150 5220 5170 5230
rect 5240 5220 5300 5240
rect 4130 5210 5160 5220
rect 2000 5200 3510 5210
rect 4110 5200 5160 5210
rect 2000 5190 3520 5200
rect 4090 5190 5160 5200
rect 2010 5180 3590 5190
rect 4080 5180 5160 5190
rect 2010 5170 3660 5180
rect 4060 5170 5160 5180
rect 2020 5160 3680 5170
rect 3750 5169 3780 5170
rect 3741 5160 3780 5169
rect 4030 5160 5160 5170
rect 2030 5150 3750 5160
rect 4020 5150 5160 5160
rect 2030 5140 3710 5150
rect 4000 5140 5160 5150
rect 2030 5130 3660 5140
rect 3990 5130 5160 5140
rect 2030 5120 3630 5130
rect 3970 5120 5160 5130
rect 2030 5110 3610 5120
rect 3960 5110 5160 5120
rect 5230 5120 5300 5220
rect 5230 5110 5290 5120
rect 2030 5100 3600 5110
rect 3940 5100 5160 5110
rect 2030 5090 3570 5100
rect 3940 5090 5170 5100
rect 2030 5080 3550 5090
rect 3920 5080 5170 5090
rect 2040 5070 3550 5080
rect 2040 5030 3560 5070
rect 3910 5060 5170 5080
rect 5220 5070 5290 5110
rect 3900 5050 4660 5060
rect 4680 5050 5170 5060
rect 3890 5040 4650 5050
rect 4700 5040 5170 5050
rect 5230 5050 5290 5070
rect 5230 5040 5280 5050
rect 3890 5030 4640 5040
rect 4720 5030 5170 5040
rect 5220 5030 5280 5040
rect 2050 5020 3560 5030
rect 3680 5020 3730 5030
rect 3840 5020 3860 5030
rect 2050 5010 3570 5020
rect 3670 5010 3770 5020
rect 3820 5010 3860 5020
rect 3880 5020 4640 5030
rect 4730 5020 5170 5030
rect 3880 5010 4630 5020
rect 2050 5000 3860 5010
rect 3870 5000 4630 5010
rect 4740 5000 5170 5020
rect 5230 5010 5280 5030
rect 5220 5000 5270 5010
rect 2060 4990 2550 5000
rect 2600 4990 4630 5000
rect 4760 4990 5170 5000
rect 2070 4980 2520 4990
rect 2620 4980 4620 4990
rect 4770 4980 5160 4990
rect 5200 4980 5270 5000
rect 2070 4970 2510 4980
rect 2630 4970 4620 4980
rect 2080 4960 2500 4970
rect 2640 4960 4620 4970
rect 4780 4970 5170 4980
rect 5200 4970 5260 4980
rect 4780 4960 5260 4970
rect 2080 4950 2490 4960
rect 2650 4950 4620 4960
rect 4790 4950 5260 4960
rect 2090 4930 2480 4950
rect 2660 4940 4620 4950
rect 2670 4930 4620 4940
rect 4800 4930 5250 4950
rect 2100 4920 2470 4930
rect 2690 4920 4620 4930
rect 2100 4910 2460 4920
rect 2700 4910 4620 4920
rect 4810 4910 5240 4930
rect 2100 4890 2450 4910
rect 2730 4900 4610 4910
rect 4820 4900 5240 4910
rect 2750 4890 4610 4900
rect 2110 4870 2450 4890
rect 2770 4880 4610 4890
rect 4830 4880 5230 4900
rect 2780 4870 4610 4880
rect 4840 4870 5220 4880
rect 2110 4850 2440 4870
rect 2790 4860 4600 4870
rect 2800 4850 4600 4860
rect 4850 4860 5220 4870
rect 4850 4850 5210 4860
rect 2120 4830 2440 4850
rect 2820 4830 4600 4850
rect 4860 4840 5200 4850
rect 2130 4820 2440 4830
rect 2830 4820 4590 4830
rect 4870 4820 5190 4840
rect 2130 4810 2450 4820
rect 2140 4790 2450 4810
rect 2150 4750 2450 4790
rect 2830 4810 3440 4820
rect 3580 4810 4590 4820
rect 4880 4810 5180 4820
rect 2830 4800 3390 4810
rect 3640 4800 4590 4810
rect 4890 4800 5170 4810
rect 2830 4790 3320 4800
rect 3660 4790 3700 4800
rect 3740 4790 4580 4800
rect 4890 4790 5160 4800
rect 2830 4770 3300 4790
rect 3760 4780 4580 4790
rect 4900 4780 5150 4790
rect 3770 4770 4580 4780
rect 4910 4770 5140 4780
rect 2830 4750 3290 4770
rect 3780 4750 4570 4770
rect 4920 4760 5120 4770
rect 4930 4750 5100 4760
rect 2150 4730 2460 4750
rect 2820 4740 3290 4750
rect 2140 4720 2460 4730
rect 2810 4730 2890 4740
rect 2910 4730 3300 4740
rect 3790 4730 4570 4750
rect 4940 4740 5080 4750
rect 4960 4730 5060 4740
rect 2810 4720 2860 4730
rect 2140 4700 2470 4720
rect 2820 4710 2850 4720
rect 2940 4710 3310 4730
rect 3800 4710 4570 4730
rect 4970 4720 5040 4730
rect 4990 4710 5030 4720
rect 2930 4700 3320 4710
rect 3800 4700 4560 4710
rect 2140 4690 2480 4700
rect 2130 4680 2480 4690
rect 2930 4690 3330 4700
rect 2930 4680 3340 4690
rect 3810 4680 4560 4700
rect 2130 4670 2490 4680
rect 2930 4670 3350 4680
rect 3810 4670 4550 4680
rect 2130 4650 2500 4670
rect 2920 4660 3370 4670
rect 3820 4660 4550 4670
rect 2920 4650 2950 4660
rect 3000 4650 3380 4660
rect 3820 4650 4540 4660
rect 2130 4630 2510 4650
rect 2920 4640 2940 4650
rect 3020 4640 3380 4650
rect 2920 4630 2930 4640
rect 3040 4630 3380 4640
rect 2130 4620 2520 4630
rect 3060 4620 3380 4630
rect 3830 4620 4520 4650
rect 2140 4600 2530 4620
rect 2140 4590 2540 4600
rect 3070 4590 3380 4620
rect 3840 4610 4510 4620
rect 3850 4600 4510 4610
rect 3860 4590 4510 4600
rect 2150 4580 2540 4590
rect 2160 4570 2550 4580
rect 2910 4570 2920 4590
rect 3080 4570 3380 4590
rect 3870 4580 4500 4590
rect 3890 4570 4400 4580
rect 4430 4570 4500 4580
rect 2170 4560 2560 4570
rect 2910 4560 2930 4570
rect 2190 4550 2610 4560
rect 2210 4540 2610 4550
rect 2910 4540 2940 4560
rect 3080 4550 3390 4570
rect 3890 4560 4380 4570
rect 4440 4560 4500 4570
rect 3910 4550 4340 4560
rect 4450 4550 4500 4560
rect 3080 4540 3400 4550
rect 3920 4540 4310 4550
rect 4450 4540 4510 4550
rect 2220 4530 2620 4540
rect 2910 4530 2950 4540
rect 2220 4520 2630 4530
rect 2910 4520 2960 4530
rect 3090 4520 3400 4540
rect 3990 4530 4290 4540
rect 4070 4520 4270 4530
rect 4460 4520 4510 4540
rect 4660 4530 4780 4540
rect 4640 4520 4800 4530
rect 2230 4510 2640 4520
rect 2920 4510 2990 4520
rect 2290 4500 2650 4510
rect 2930 4500 3000 4510
rect 3090 4500 3390 4520
rect 4090 4510 4240 4520
rect 4460 4510 4520 4520
rect 4630 4510 4820 4520
rect 4120 4500 4200 4510
rect 4470 4500 4550 4510
rect 4610 4500 4830 4510
rect 2320 4490 2660 4500
rect 2930 4490 3020 4500
rect 3090 4490 3380 4500
rect 3440 4490 3500 4500
rect 4470 4490 4570 4500
rect 4580 4490 4840 4500
rect 2340 4480 2660 4490
rect 2360 4470 2670 4480
rect 2940 4470 3030 4490
rect 2360 4460 2680 4470
rect 2960 4460 3020 4470
rect 3090 4460 3370 4490
rect 3440 4460 3510 4490
rect 4480 4480 4840 4490
rect 4490 4470 4840 4480
rect 4510 4460 4840 4470
rect 2370 4450 2690 4460
rect 3090 4450 3380 4460
rect 3440 4450 3500 4460
rect 4530 4450 4840 4460
rect 2370 4440 2700 4450
rect 2360 4430 2700 4440
rect 3080 4430 3380 4450
rect 3430 4440 3490 4450
rect 4550 4440 4830 4450
rect 3430 4430 3480 4440
rect 4560 4430 4680 4440
rect 4750 4430 4830 4440
rect 2360 4420 2710 4430
rect 2360 4400 2720 4420
rect 3070 4410 3380 4430
rect 3420 4420 3480 4430
rect 3420 4410 3460 4420
rect 4760 4410 4830 4430
rect 2360 4390 2730 4400
rect 3060 4390 3390 4410
rect 4760 4400 4820 4410
rect 4760 4390 4810 4400
rect 2360 4380 2740 4390
rect 3070 4380 3400 4390
rect 2370 4370 2750 4380
rect 3080 4370 3400 4380
rect 2370 4360 2760 4370
rect 3090 4360 3400 4370
rect 2370 4350 2770 4360
rect 3100 4350 3410 4360
rect 3460 4350 3480 4360
rect 2380 4340 2780 4350
rect 3100 4340 3420 4350
rect 3450 4340 3480 4350
rect 2380 4330 2800 4340
rect 3110 4330 3430 4340
rect 3440 4330 3480 4340
rect 2400 4320 2810 4330
rect 3110 4320 3460 4330
rect 2410 4310 2830 4320
rect 2430 4300 2840 4310
rect 2460 4290 2850 4300
rect 2470 4280 2860 4290
rect 3120 4280 3450 4320
rect 2470 4270 2870 4280
rect 3110 4270 3450 4280
rect 2460 4260 2890 4270
rect 3100 4260 3450 4270
rect 4970 4260 4990 4270
rect 2450 4250 2910 4260
rect 3080 4250 3510 4260
rect 4930 4250 4990 4260
rect 2450 4240 2940 4250
rect 3060 4240 3520 4250
rect 4910 4240 4990 4250
rect 2450 4230 2980 4240
rect 3040 4230 3520 4240
rect 2450 4220 3520 4230
rect 4890 4220 4990 4240
rect 2460 4210 3520 4220
rect 4600 4210 4650 4220
rect 4820 4210 4990 4220
rect 2460 4200 3530 4210
rect 4560 4200 4670 4210
rect 4720 4200 4980 4210
rect 2470 4190 3530 4200
rect 4510 4190 4900 4200
rect 2470 4180 3470 4190
rect 3480 4180 3530 4190
rect 4460 4180 4880 4190
rect 2480 4170 3470 4180
rect 2490 4160 3470 4170
rect 3500 4160 3520 4180
rect 4370 4170 4830 4180
rect 4350 4160 4610 4170
rect 4640 4160 4820 4170
rect 2500 4150 3480 4160
rect 2510 4140 3480 4150
rect 4340 4150 4570 4160
rect 4340 4140 4540 4150
rect 2510 4130 3490 4140
rect 4330 4130 4530 4140
rect 2520 4120 3500 4130
rect 2540 4110 3500 4120
rect 4330 4120 4490 4130
rect 4330 4110 4450 4120
rect 2550 4100 3510 4110
rect 2570 4090 3520 4100
rect 2580 4080 3530 4090
rect 2590 4070 3540 4080
rect 2600 4060 3550 4070
rect 2610 4050 3560 4060
rect 2620 4040 3560 4050
rect 4810 4040 4880 4050
rect 2630 4030 3570 4040
rect 4770 4030 4880 4040
rect 2640 4020 3580 4030
rect 4720 4020 4890 4030
rect 2660 4010 3590 4020
rect 4650 4010 4880 4020
rect 2700 4000 3600 4010
rect 4630 4000 4880 4010
rect 2720 3990 2760 4000
rect 2800 3990 3610 4000
rect 4610 3990 4870 4000
rect 2810 3980 3610 3990
rect 4580 3980 4860 3990
rect 2810 3970 3620 3980
rect 4570 3970 4840 3980
rect 2820 3960 3630 3970
rect 4580 3960 4810 3970
rect 2820 3950 3650 3960
rect 4610 3950 4650 3960
rect 2830 3940 3670 3950
rect 2850 3930 3720 3940
rect 2880 3920 3730 3930
rect 2930 3910 3740 3920
rect 2950 3900 3760 3910
rect 2950 3890 3780 3900
rect 2950 3880 3800 3890
rect 2950 3870 3830 3880
rect 2950 3860 3880 3870
rect 2950 3850 3900 3860
rect 2950 3840 3950 3850
rect 2950 3830 4010 3840
rect 2950 3820 4030 3830
rect 2950 3810 4040 3820
rect 2950 3800 4080 3810
rect 2950 3780 4090 3800
rect 4490 3780 4550 3790
rect 2950 3770 4100 3780
rect 4470 3770 4540 3780
rect 2950 3760 4110 3770
rect 4170 3760 4180 3770
rect 4440 3760 4530 3770
rect 2950 3750 4120 3760
rect 4140 3750 4230 3760
rect 4250 3750 4290 3760
rect 4360 3750 4520 3760
rect 2950 3740 4510 3750
rect 2950 3730 4490 3740
rect 2950 3720 4480 3730
rect 2940 3710 4460 3720
rect 2940 3700 4440 3710
rect 2940 3690 4430 3700
rect 2940 3680 4420 3690
rect 2940 3670 4410 3680
rect 2940 3660 4400 3670
rect 2940 3650 4390 3660
rect 4970 3650 4990 3660
rect 2940 3640 4380 3650
rect 4940 3640 5000 3650
rect 2930 3630 4380 3640
rect 4920 3630 4980 3640
rect 2930 3620 4370 3630
rect 4910 3620 4970 3630
rect 2930 3610 4360 3620
rect 4900 3610 4960 3620
rect 2920 3600 4350 3610
rect 4910 3600 4940 3610
rect 2920 3590 4340 3600
rect 2920 3580 4330 3590
rect 2910 3570 4330 3580
rect 2910 3560 3320 3570
rect 3330 3560 4320 3570
rect 2900 3550 3310 3560
rect 3340 3550 4310 3560
rect 2890 3540 3310 3550
rect 3410 3540 4300 3550
rect 2890 3530 3300 3540
rect 3420 3530 4290 3540
rect 2880 3520 3300 3530
rect 3430 3520 4280 3530
rect 2880 3510 3290 3520
rect 3450 3510 4270 3520
rect 2870 3500 3290 3510
rect 3470 3500 4260 3510
rect 2870 3490 3260 3500
rect 3490 3490 4250 3500
rect 2860 3480 3250 3490
rect 3500 3480 4240 3490
rect 2850 3470 3240 3480
rect 3520 3470 4230 3480
rect 2840 3450 3240 3470
rect 3530 3460 4220 3470
rect 3540 3450 4200 3460
rect 2830 3440 3240 3450
rect 3550 3440 4190 3450
rect 2600 3430 2670 3440
rect 2840 3430 2860 3440
rect 2910 3430 3250 3440
rect 3550 3430 4180 3440
rect 2580 3420 2700 3430
rect 2910 3420 3290 3430
rect 3550 3420 4160 3430
rect 2560 3410 2710 3420
rect 2920 3410 3300 3420
rect 3560 3410 4150 3420
rect 2550 3400 2700 3410
rect 2960 3400 3290 3410
rect 3570 3400 4140 3410
rect 2530 3390 2700 3400
rect 3000 3390 3260 3400
rect 3600 3390 4130 3400
rect 2520 3380 2690 3390
rect 3010 3380 3250 3390
rect 3610 3380 4120 3390
rect 2500 3370 2690 3380
rect 3040 3370 3250 3380
rect 3630 3370 4110 3380
rect 2470 3360 2690 3370
rect 3050 3360 3240 3370
rect 2460 3350 2690 3360
rect 3060 3350 3240 3360
rect 3650 3360 4100 3370
rect 3650 3350 4090 3360
rect 2430 3340 2690 3350
rect 3090 3340 3230 3350
rect 2410 3330 2690 3340
rect 3100 3330 3230 3340
rect 3660 3340 4070 3350
rect 3660 3330 4060 3340
rect 2400 3320 2700 3330
rect 2380 3310 2700 3320
rect 3100 3320 3220 3330
rect 3100 3310 3180 3320
rect 3670 3310 4050 3330
rect 2360 3300 2700 3310
rect 3110 3300 3170 3310
rect 3670 3300 4040 3310
rect 2340 3290 2710 3300
rect 3140 3290 3150 3300
rect 3660 3290 4030 3300
rect 2320 3280 2720 3290
rect 3650 3280 4020 3290
rect 2300 3270 2730 3280
rect 3640 3270 4010 3280
rect 2280 3260 2740 3270
rect 3630 3260 4000 3270
rect 2250 3250 2740 3260
rect 3510 3250 3520 3260
rect 3600 3250 4000 3260
rect 2230 3240 2750 3250
rect 3500 3240 3530 3250
rect 2210 3230 2760 3240
rect 3510 3230 3530 3240
rect 3580 3240 3990 3250
rect 2190 3220 2760 3230
rect 3580 3220 3980 3240
rect 2170 3210 2770 3220
rect 3580 3210 3970 3220
rect 2140 3200 2780 3210
rect 3510 3200 3560 3210
rect 3570 3200 3970 3210
rect 2120 3190 2790 3200
rect 3510 3190 3960 3200
rect 2090 3180 2800 3190
rect 3510 3180 3950 3190
rect 2050 3170 2800 3180
rect 3550 3170 3950 3180
rect 2020 3160 2810 3170
rect 3550 3160 3940 3170
rect 4870 3160 4900 3170
rect 1990 3150 2820 3160
rect 3540 3150 3930 3160
rect 4870 3150 4880 3160
rect 1960 3140 2840 3150
rect 1930 3130 2850 3140
rect 3540 3130 3920 3150
rect 1890 3120 2860 3130
rect 3540 3120 3910 3130
rect 1840 3110 2870 3120
rect 3550 3110 3900 3120
rect 1800 3100 2890 3110
rect 1750 3090 2900 3100
rect 3550 3090 3890 3110
rect 1720 3080 2910 3090
rect 3550 3080 3880 3090
rect 1690 3070 2920 3080
rect 1650 3060 2920 3070
rect 3550 3070 3870 3080
rect 3550 3060 3860 3070
rect 1620 3050 2930 3060
rect 3560 3050 3860 3060
rect 1590 3040 2950 3050
rect 3570 3040 3860 3050
rect 1540 3030 2960 3040
rect 1510 3020 2980 3030
rect 3370 3020 3410 3030
rect 3580 3020 3610 3040
rect 3630 3020 3850 3040
rect 1460 3010 3000 3020
rect 1400 3000 3010 3010
rect 3360 3000 3420 3020
rect 3560 3010 3840 3020
rect 1370 2990 3030 3000
rect 3350 2990 3420 3000
rect 3550 3000 3840 3010
rect 1320 2980 3040 2990
rect 3360 2980 3410 2990
rect 1270 2970 3050 2980
rect 3380 2970 3400 2980
rect 3550 2970 3830 3000
rect 1240 2960 3070 2970
rect 3540 2960 3830 2970
rect 1190 2950 3090 2960
rect 3530 2950 3830 2960
rect 1160 2940 3100 2950
rect 3520 2940 3820 2950
rect 1130 2930 3130 2940
rect 3510 2930 3820 2940
rect 1100 2920 3160 2930
rect 3320 2920 3340 2930
rect 3500 2920 3820 2930
rect 1080 2910 3170 2920
rect 1070 2900 3180 2910
rect 3310 2900 3360 2920
rect 3490 2910 3830 2920
rect 3470 2900 3830 2910
rect 1050 2890 3200 2900
rect 3250 2890 3360 2900
rect 3440 2890 3820 2900
rect 1040 2880 3370 2890
rect 3420 2880 3820 2890
rect 1030 2870 3370 2880
rect 1010 2860 3370 2870
rect 1000 2850 3370 2860
rect 3410 2870 3820 2880
rect 990 2840 3360 2850
rect 970 2830 3360 2840
rect 960 2820 3370 2830
rect 960 2810 3380 2820
rect 3410 2810 3830 2870
rect 950 2800 3830 2810
rect 940 2790 3830 2800
rect 930 2780 3830 2790
rect 920 2770 3440 2780
rect 3470 2770 3830 2780
rect 910 2760 3830 2770
rect 910 2750 3840 2760
rect 900 2730 3840 2750
rect 5190 2730 5240 2740
rect 890 2720 3840 2730
rect 5180 2720 5270 2730
rect 880 2700 3840 2720
rect 5170 2710 5280 2720
rect 5160 2700 5300 2710
rect 870 2690 3840 2700
rect 5150 2690 5310 2700
rect 860 2680 3830 2690
rect 5140 2680 5330 2690
rect 850 2660 3830 2680
rect 5120 2670 5340 2680
rect 5110 2660 5350 2670
rect 840 2640 3830 2660
rect 5090 2650 5370 2660
rect 5070 2640 5390 2650
rect 830 2630 3830 2640
rect 5060 2630 5400 2640
rect 820 2620 3830 2630
rect 5040 2620 5420 2630
rect 820 2610 3820 2620
rect 5030 2610 5440 2620
rect 810 2590 3820 2610
rect 5020 2600 5450 2610
rect 5010 2590 5470 2600
rect 800 2580 3820 2590
rect 5000 2580 5490 2590
rect 790 2560 3810 2580
rect 4990 2570 5510 2580
rect 4990 2560 5530 2570
rect 780 2540 3810 2560
rect 4980 2550 5550 2560
rect 4970 2540 5570 2550
rect 770 2510 3810 2540
rect 4960 2530 5590 2540
rect 4950 2520 5600 2530
rect 760 2480 3800 2510
rect 4940 2500 5610 2520
rect 4940 2490 5620 2500
rect 750 2460 3790 2480
rect 4930 2470 5630 2490
rect 740 2440 3790 2460
rect 4920 2460 5640 2470
rect 4920 2450 5650 2460
rect 4880 2440 4890 2450
rect 4910 2440 5650 2450
rect 740 2420 3780 2440
rect 4870 2430 5660 2440
rect 4860 2420 5670 2430
rect 730 2400 3780 2420
rect 4850 2410 5670 2420
rect 4850 2400 5680 2410
rect 730 2380 3770 2400
rect 4850 2390 5690 2400
rect 720 2370 3770 2380
rect 4840 2380 5690 2390
rect 4840 2370 5700 2380
rect 720 2350 3760 2370
rect 4830 2360 5710 2370
rect 710 2330 3760 2350
rect 4820 2350 5710 2360
rect 4820 2340 5720 2350
rect 4810 2330 5720 2340
rect 710 2310 3750 2330
rect 4810 2320 5730 2330
rect 4800 2310 5740 2320
rect 700 2300 3750 2310
rect 4790 2300 5740 2310
rect 700 2290 3740 2300
rect 4780 2290 5750 2300
rect 690 2280 3740 2290
rect 4770 2280 5760 2290
rect 690 2260 3730 2280
rect 4760 2270 5760 2280
rect 4760 2260 5770 2270
rect 680 2250 3730 2260
rect 4750 2250 5770 2260
rect 680 2230 3720 2250
rect 4740 2230 5780 2250
rect 670 2220 3710 2230
rect 670 2200 3700 2220
rect 4730 2210 5790 2230
rect 4720 2200 5790 2210
rect 670 2190 3690 2200
rect 4710 2190 5790 2200
rect 660 2170 3680 2190
rect 4700 2180 5800 2190
rect 4690 2170 5800 2180
rect 660 2150 3670 2170
rect 4680 2160 5800 2170
rect 4670 2150 5810 2160
rect 660 2140 3660 2150
rect 4660 2140 5810 2150
rect 650 2130 3660 2140
rect 4650 2130 5810 2140
rect 650 2110 3650 2130
rect 4640 2110 5820 2130
rect 650 2100 3640 2110
rect 4620 2100 5820 2110
rect 650 2080 3630 2100
rect 4610 2090 5820 2100
rect 4600 2080 5820 2090
rect 650 2070 3620 2080
rect 4580 2070 5820 2080
rect 640 2040 3610 2070
rect 4570 2060 5820 2070
rect 4550 2050 5830 2060
rect 640 2020 3600 2040
rect 4540 2030 5830 2050
rect 5990 2040 6000 2220
rect 4530 2020 5830 2030
rect 640 2010 3590 2020
rect 4520 2010 5830 2020
rect 630 2000 3590 2010
rect 4510 2000 5830 2010
rect 630 1980 3580 2000
rect 4500 1990 5840 2000
rect 4490 1980 5840 1990
rect 630 1970 3570 1980
rect 4480 1970 5840 1980
rect 630 1950 3560 1970
rect 4470 1960 5840 1970
rect 4460 1950 5840 1960
rect 630 1930 3550 1950
rect 4450 1940 5840 1950
rect 630 1920 3540 1930
rect 4450 1920 5850 1940
rect 620 1900 3530 1920
rect 4440 1900 5850 1920
rect 620 1890 3520 1900
rect 4430 1890 5850 1900
rect 620 1870 3510 1890
rect 4430 1880 5860 1890
rect 620 1860 3500 1870
rect 4420 1860 5860 1880
rect 620 1840 3490 1860
rect 4410 1850 5870 1860
rect 620 1820 3480 1840
rect 4400 1830 5870 1850
rect 4390 1820 5870 1830
rect 620 1800 3470 1820
rect 4380 1810 5870 1820
rect 4370 1800 5880 1810
rect 620 1780 3460 1800
rect 4360 1790 5880 1800
rect 4350 1780 5880 1790
rect 620 1760 3450 1780
rect 4340 1760 5880 1780
rect 620 1740 3440 1760
rect 4330 1750 5880 1760
rect 620 1720 3430 1740
rect 4320 1730 5890 1750
rect 4310 1720 5890 1730
rect 620 1700 3420 1720
rect 4300 1700 5890 1720
rect 620 1680 3410 1700
rect 4290 1690 5890 1700
rect 4290 1680 5900 1690
rect 620 1660 3400 1680
rect 4280 1670 5900 1680
rect 620 1640 3390 1660
rect 4270 1650 5900 1670
rect 620 1620 3380 1640
rect 4270 1630 5910 1650
rect 4260 1620 4400 1630
rect 4450 1620 5910 1630
rect 620 1600 3370 1620
rect 4260 1610 4390 1620
rect 4460 1610 5910 1620
rect 4250 1600 4380 1610
rect 4470 1600 5910 1610
rect 620 1580 3360 1600
rect 4250 1590 4370 1600
rect 4490 1590 5910 1600
rect 4240 1580 4360 1590
rect 4500 1580 5910 1590
rect 620 1560 3350 1580
rect 4240 1570 4350 1580
rect 4510 1570 5920 1580
rect 4240 1560 4340 1570
rect 4530 1560 5920 1570
rect 620 1540 3340 1560
rect 4240 1550 4330 1560
rect 4540 1550 5920 1560
rect 4230 1540 4320 1550
rect 4550 1540 5920 1550
rect 620 1520 3330 1540
rect 4230 1530 4310 1540
rect 4560 1530 5920 1540
rect 4220 1520 4300 1530
rect 4570 1520 5930 1530
rect 620 1500 3320 1520
rect 4220 1510 4290 1520
rect 4580 1510 5930 1520
rect 4220 1500 4280 1510
rect 4590 1500 5930 1510
rect 630 1480 3310 1500
rect 4210 1490 4260 1500
rect 4600 1490 5930 1500
rect 4210 1480 4250 1490
rect 4610 1480 5940 1490
rect 630 1460 3300 1480
rect 4210 1470 4230 1480
rect 4620 1470 5940 1480
rect 4630 1460 5940 1470
rect 630 1440 3290 1460
rect 4640 1440 5940 1460
rect 630 1410 3280 1440
rect 4650 1430 5940 1440
rect 4660 1420 5940 1430
rect 4680 1410 5940 1420
rect 640 1390 3270 1410
rect 4690 1400 5950 1410
rect 4700 1390 5950 1400
rect 640 1370 3260 1390
rect 4710 1380 5950 1390
rect 4720 1370 5950 1380
rect 640 1360 3250 1370
rect 4730 1360 5950 1370
rect 650 1350 3250 1360
rect 650 1330 3240 1350
rect 4740 1340 5960 1360
rect 4750 1330 5960 1340
rect 650 1320 3230 1330
rect 4760 1320 5960 1330
rect 650 1300 3220 1320
rect 4770 1310 5960 1320
rect 4780 1300 5960 1310
rect 650 1290 3210 1300
rect 4780 1290 5970 1300
rect 650 1270 3200 1290
rect 4790 1280 5970 1290
rect 660 1250 3190 1270
rect 4800 1260 5970 1280
rect 660 1230 3180 1250
rect 4810 1240 5970 1260
rect 4120 1230 4170 1240
rect 670 1210 3170 1230
rect 4110 1220 4200 1230
rect 4820 1220 5980 1240
rect 4100 1210 4210 1220
rect 670 1200 3160 1210
rect 4100 1200 4230 1210
rect 670 1190 3150 1200
rect 680 1180 3150 1190
rect 4090 1190 4240 1200
rect 4830 1190 5980 1220
rect 4090 1180 4250 1190
rect 680 1160 3140 1180
rect 4080 1170 4270 1180
rect 4830 1170 5990 1190
rect 4080 1160 4290 1170
rect 680 1150 3130 1160
rect 4080 1150 4300 1160
rect 4820 1150 5990 1170
rect 690 1130 3120 1150
rect 4080 1140 4310 1150
rect 4080 1130 4330 1140
rect 4810 1130 6000 1150
rect 690 1110 3110 1130
rect 4070 1120 4340 1130
rect 4800 1120 6000 1130
rect 4070 1110 4360 1120
rect 4790 1110 6000 1120
rect 700 1100 3100 1110
rect 4070 1100 4370 1110
rect 700 1080 3090 1100
rect 4060 1090 4390 1100
rect 4780 1090 6000 1110
rect 4060 1080 4410 1090
rect 4770 1080 6000 1090
rect 700 1060 3080 1080
rect 4050 1070 4430 1080
rect 4050 1060 4440 1070
rect 4760 1060 6000 1080
rect 710 1050 3070 1060
rect 4040 1050 4460 1060
rect 4750 1050 6000 1060
rect 710 1030 3060 1050
rect 4040 1040 4480 1050
rect 4740 1040 6000 1050
rect 4030 1030 4490 1040
rect 4730 1030 6000 1040
rect 710 1010 3050 1030
rect 4030 1020 4500 1030
rect 4720 1020 6000 1030
rect 4030 1010 4520 1020
rect 4710 1010 6000 1020
rect 710 1000 3040 1010
rect 4020 1000 4530 1010
rect 4700 1000 6000 1010
rect 710 980 3030 1000
rect 4020 990 4540 1000
rect 4690 990 6000 1000
rect 4020 980 4550 990
rect 4680 980 6000 990
rect 720 970 3020 980
rect 4020 970 4570 980
rect 4660 970 6000 980
rect 720 950 3010 970
rect 4010 960 4590 970
rect 4650 960 6000 970
rect 4010 950 4600 960
rect 4640 950 6000 960
rect 720 940 3000 950
rect 720 920 2990 940
rect 4000 930 4600 950
rect 4620 940 6000 950
rect 4610 930 6000 940
rect 4000 920 4590 930
rect 720 910 2980 920
rect 3990 910 4580 920
rect 4620 910 6000 930
rect 720 890 2970 910
rect 3990 900 4560 910
rect 4630 900 6000 910
rect 3990 890 4550 900
rect 4650 890 6000 900
rect 720 880 2960 890
rect 3980 880 4530 890
rect 4670 880 6000 890
rect 720 870 2950 880
rect 3980 870 4520 880
rect 4680 870 6000 880
rect 720 850 2940 870
rect 3980 860 4510 870
rect 4690 860 6000 870
rect 3970 850 4490 860
rect 4700 850 6000 860
rect 720 830 2930 850
rect 3970 840 4480 850
rect 4710 840 6000 850
rect 3960 830 4470 840
rect 4720 830 6000 840
rect 720 820 2920 830
rect 3960 820 4450 830
rect 4730 820 6000 830
rect 720 800 2910 820
rect 3960 810 4440 820
rect 4750 810 6000 820
rect 3950 800 4420 810
rect 4760 800 6000 810
rect 730 790 2900 800
rect 3950 790 4410 800
rect 4770 790 6000 800
rect 730 780 2890 790
rect 3940 780 4400 790
rect 730 770 2880 780
rect 3940 770 4380 780
rect 4780 770 6000 790
rect 730 750 2870 770
rect 3940 760 4370 770
rect 4790 760 6000 770
rect 3930 750 4360 760
rect 4800 750 6000 760
rect 730 730 2860 750
rect 3920 740 4340 750
rect 4810 740 6000 750
rect 3920 730 4320 740
rect 4820 730 6000 740
rect 730 720 2850 730
rect 3920 720 4310 730
rect 4830 720 6000 730
rect 720 710 2840 720
rect 3920 710 3940 720
rect 3980 710 4290 720
rect 4840 710 6000 720
rect 720 690 2830 710
rect 3990 700 4280 710
rect 4850 700 6000 710
rect 4010 690 4260 700
rect 4860 690 6000 700
rect 720 680 2820 690
rect 4020 680 4250 690
rect 4870 680 6000 690
rect 720 670 2810 680
rect 4030 670 4230 680
rect 720 660 2800 670
rect 4040 660 4220 670
rect 4880 660 6000 680
rect 720 640 2790 660
rect 4050 650 4200 660
rect 4060 640 4190 650
rect 720 630 2780 640
rect 4060 630 4180 640
rect 720 610 2770 630
rect 4070 620 4170 630
rect 4080 610 4160 620
rect 720 600 2760 610
rect 4090 600 4140 610
rect 730 590 2750 600
rect 4100 590 4130 600
rect 730 580 2740 590
rect 730 570 2730 580
rect 730 560 1900 570
rect 2180 560 2720 570
rect 730 550 1790 560
rect 2240 550 2710 560
rect 4890 550 6000 660
rect 730 540 1730 550
rect 2290 540 2700 550
rect 4880 540 6000 550
rect 730 530 1690 540
rect 2320 530 2690 540
rect 740 520 1660 530
rect 2350 520 2680 530
rect 4870 520 6000 540
rect 740 510 1630 520
rect 2380 510 2670 520
rect 4110 510 4130 520
rect 4860 510 6000 520
rect 730 500 1590 510
rect 2400 500 2670 510
rect 730 490 1550 500
rect 2420 490 2660 500
rect 4090 490 4140 510
rect 4850 500 6000 510
rect 4840 490 6000 500
rect 730 480 1520 490
rect 2430 480 2640 490
rect 4080 480 4140 490
rect 4830 480 6000 490
rect 730 470 1500 480
rect 2440 470 2630 480
rect 4070 470 4140 480
rect 4820 470 6000 480
rect 730 460 1480 470
rect 730 450 1460 460
rect 2450 450 2620 470
rect 4060 460 4130 470
rect 4810 460 6000 470
rect 4060 450 4120 460
rect 4800 450 6000 460
rect 730 440 1450 450
rect 2460 440 2610 450
rect 4050 440 4120 450
rect 4780 440 6000 450
rect 730 430 1430 440
rect 2470 430 2600 440
rect 4050 430 4100 440
rect 4160 430 4170 440
rect 4770 430 6000 440
rect 730 420 1420 430
rect 2470 420 2590 430
rect 4040 420 4090 430
rect 4150 420 4180 430
rect 4760 420 6000 430
rect 730 410 1410 420
rect 2470 410 2580 420
rect 4030 410 4090 420
rect 4160 410 4190 420
rect 4740 410 6000 420
rect 730 400 1400 410
rect 2480 400 2570 410
rect 730 380 1390 400
rect 2480 390 2560 400
rect 4020 390 4080 410
rect 4160 400 4200 410
rect 4730 400 6000 410
rect 4170 390 4200 400
rect 4720 390 6000 400
rect 2480 380 2540 390
rect 4010 380 4070 390
rect 4710 380 6000 390
rect 740 370 1380 380
rect 2500 370 2510 380
rect 4000 370 4060 380
rect 4700 370 6000 380
rect 740 340 1370 370
rect 3990 360 4050 370
rect 4690 360 6000 370
rect 3980 350 4040 360
rect 4670 350 6000 360
rect 3970 340 4030 350
rect 4660 340 6000 350
rect 740 330 1360 340
rect 3960 330 4030 340
rect 4640 330 6000 340
rect 730 320 1350 330
rect 3950 320 4010 330
rect 4630 320 6000 330
rect 740 310 1350 320
rect 3940 310 4010 320
rect 4280 310 4290 320
rect 4620 310 6000 320
rect 740 300 1340 310
rect 3940 300 4000 310
rect 4280 300 4300 310
rect 4600 300 6000 310
rect 740 280 1330 300
rect 3930 290 3990 300
rect 4290 290 4300 300
rect 4580 290 6000 300
rect 3920 280 3980 290
rect 4570 280 6000 290
rect 740 250 1320 280
rect 3910 270 3970 280
rect 4550 270 6000 280
rect 3900 260 3960 270
rect 4320 260 4340 270
rect 4540 260 6000 270
rect 3890 250 3950 260
rect 4330 250 4350 260
rect 4520 250 6000 260
rect 740 220 1310 250
rect 3880 240 3940 250
rect 4340 240 4360 250
rect 4500 240 6000 250
rect 3870 230 3930 240
rect 4350 230 4380 240
rect 4490 230 6000 240
rect 3860 220 3920 230
rect 4360 220 4400 230
rect 4470 220 6000 230
rect 740 200 1300 220
rect 3720 210 3790 220
rect 3850 210 3910 220
rect 4370 210 4420 220
rect 4440 210 4570 220
rect 3720 200 3810 210
rect 3840 200 3900 210
rect 4380 200 4550 210
rect 740 180 1290 200
rect 3710 190 3890 200
rect 4390 190 4540 200
rect 4610 190 6000 220
rect 3720 180 3880 190
rect 4400 180 4520 190
rect 750 160 1290 180
rect 3750 170 3870 180
rect 4400 170 4500 180
rect 3770 160 3870 170
rect 4410 160 4490 170
rect 4600 160 6000 190
rect 760 150 1280 160
rect 3780 150 3860 160
rect 4420 150 4470 160
rect 780 140 1280 150
rect 3790 140 3850 150
rect 4430 140 4450 150
rect 790 130 1280 140
rect 3800 130 3830 140
rect 4590 130 6000 160
rect 810 120 1280 130
rect 830 110 1280 120
rect 4580 120 5970 130
rect 4580 110 5960 120
rect 850 100 1280 110
rect 4560 100 5930 110
rect 870 90 1280 100
rect 4550 90 5900 100
rect 880 80 1280 90
rect 4540 80 5880 90
rect 910 70 1280 80
rect 4520 70 5820 80
rect 950 60 1270 70
rect 4510 60 5760 70
rect 1000 50 1220 60
rect 1240 50 1270 60
rect 3660 50 3710 60
rect 4500 50 5730 60
rect 3650 40 3730 50
rect 4480 40 5700 50
rect 3640 30 3750 40
rect 4470 30 5690 40
rect 3640 20 3760 30
rect 4460 20 5670 30
rect 3630 10 3780 20
rect 4450 10 5660 20
rect 3630 0 3800 10
rect 4440 0 5660 10
<< end >>
