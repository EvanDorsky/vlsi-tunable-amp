magic
tech scmos
timestamp 1259953556
<< electrodecontact >>
rect 20 4090 24 4094
rect 38 4090 42 4094
rect 64 4089 68 4093
rect 70 4089 74 4093
rect 76 4089 80 4093
rect 82 4089 86 4093
rect 89 4089 93 4093
rect 95 4089 99 4093
rect 20 4084 24 4088
rect 38 4084 42 4088
rect 64 4083 68 4087
rect 70 4083 74 4087
rect 76 4083 80 4087
rect 82 4083 86 4087
rect 89 4083 93 4087
rect 95 4083 99 4087
rect 20 4078 24 4082
rect 38 4078 42 4082
rect 64 4077 68 4081
rect 70 4077 74 4081
rect 76 4077 80 4081
rect 82 4077 86 4081
rect 89 4077 93 4081
rect 95 4077 99 4081
rect 20 4072 24 4076
rect 38 4072 42 4076
rect 64 4071 68 4075
rect 70 4071 74 4075
rect 76 4071 80 4075
rect 82 4071 86 4075
rect 89 4071 93 4075
rect 95 4071 99 4075
rect 20 4066 24 4070
rect 38 4066 42 4070
rect 64 4065 68 4069
rect 70 4065 74 4069
rect 76 4065 80 4069
rect 82 4065 86 4069
rect 89 4065 93 4069
rect 95 4065 99 4069
rect 112 4090 116 4094
rect 125 4090 129 4094
rect 112 4084 116 4088
rect 125 4084 129 4088
rect 112 4078 116 4082
rect 125 4078 129 4082
rect 112 4072 116 4076
rect 125 4072 129 4076
rect 112 4066 116 4070
rect 125 4066 129 4070
rect 20 4060 24 4064
rect 38 4060 42 4064
rect 112 4060 116 4064
rect 125 4060 129 4064
rect 20 4054 24 4058
rect 38 4054 42 4058
rect 53 4056 57 4060
rect 112 4054 116 4058
rect 125 4054 129 4058
rect 53 4046 57 4050
rect 53 4008 57 4012
rect 20 4000 24 4004
rect 38 4000 42 4004
rect 53 3998 57 4002
rect 112 4000 116 4004
rect 125 4000 129 4004
rect 20 3994 24 3998
rect 38 3994 42 3998
rect 112 3994 116 3998
rect 125 3994 129 3998
rect 20 3988 24 3992
rect 38 3988 42 3992
rect 64 3989 68 3993
rect 70 3989 74 3993
rect 76 3989 80 3993
rect 82 3989 86 3993
rect 89 3989 93 3993
rect 95 3989 99 3993
rect 20 3982 24 3986
rect 38 3982 42 3986
rect 64 3983 68 3987
rect 70 3983 74 3987
rect 76 3983 80 3987
rect 82 3983 86 3987
rect 89 3983 93 3987
rect 95 3983 99 3987
rect 20 3976 24 3980
rect 38 3976 42 3980
rect 64 3977 68 3981
rect 70 3977 74 3981
rect 76 3977 80 3981
rect 82 3977 86 3981
rect 89 3977 93 3981
rect 95 3977 99 3981
rect 20 3970 24 3974
rect 38 3970 42 3974
rect 64 3971 68 3975
rect 70 3971 74 3975
rect 76 3971 80 3975
rect 82 3971 86 3975
rect 89 3971 93 3975
rect 95 3971 99 3975
rect 20 3964 24 3968
rect 38 3964 42 3968
rect 64 3965 68 3969
rect 70 3965 74 3969
rect 76 3965 80 3969
rect 82 3965 86 3969
rect 89 3965 93 3969
rect 95 3965 99 3969
rect 112 3988 116 3992
rect 125 3988 129 3992
rect 112 3982 116 3986
rect 125 3982 129 3986
rect 112 3976 116 3980
rect 125 3976 129 3980
rect 112 3970 116 3974
rect 125 3970 129 3974
rect 112 3964 116 3968
rect 125 3964 129 3968
rect 20 3616 24 3620
rect 38 3616 42 3620
rect 64 3615 68 3619
rect 70 3615 74 3619
rect 76 3615 80 3619
rect 82 3615 86 3619
rect 89 3615 93 3619
rect 95 3615 99 3619
rect 20 3610 24 3614
rect 38 3610 42 3614
rect 64 3609 68 3613
rect 70 3609 74 3613
rect 76 3609 80 3613
rect 82 3609 86 3613
rect 89 3609 93 3613
rect 95 3609 99 3613
rect 20 3604 24 3608
rect 38 3604 42 3608
rect 64 3603 68 3607
rect 70 3603 74 3607
rect 76 3603 80 3607
rect 82 3603 86 3607
rect 89 3603 93 3607
rect 95 3603 99 3607
rect 20 3598 24 3602
rect 38 3598 42 3602
rect 64 3597 68 3601
rect 70 3597 74 3601
rect 76 3597 80 3601
rect 82 3597 86 3601
rect 89 3597 93 3601
rect 95 3597 99 3601
rect 20 3592 24 3596
rect 38 3592 42 3596
rect 64 3591 68 3595
rect 70 3591 74 3595
rect 76 3591 80 3595
rect 82 3591 86 3595
rect 89 3591 93 3595
rect 95 3591 99 3595
rect 112 3616 116 3620
rect 125 3616 129 3620
rect 112 3610 116 3614
rect 125 3610 129 3614
rect 112 3604 116 3608
rect 125 3604 129 3608
rect 112 3598 116 3602
rect 125 3598 129 3602
rect 112 3592 116 3596
rect 125 3592 129 3596
rect 20 3586 24 3590
rect 38 3586 42 3590
rect 112 3586 116 3590
rect 125 3586 129 3590
rect 20 3580 24 3584
rect 38 3580 42 3584
rect 53 3582 57 3586
rect 112 3580 116 3584
rect 125 3580 129 3584
rect 53 3572 57 3576
rect 53 3534 57 3538
rect 20 3526 24 3530
rect 38 3526 42 3530
rect 53 3524 57 3528
rect 112 3526 116 3530
rect 125 3526 129 3530
rect 20 3520 24 3524
rect 38 3520 42 3524
rect 112 3520 116 3524
rect 125 3520 129 3524
rect 20 3514 24 3518
rect 38 3514 42 3518
rect 64 3515 68 3519
rect 70 3515 74 3519
rect 76 3515 80 3519
rect 82 3515 86 3519
rect 89 3515 93 3519
rect 95 3515 99 3519
rect 20 3508 24 3512
rect 38 3508 42 3512
rect 64 3509 68 3513
rect 70 3509 74 3513
rect 76 3509 80 3513
rect 82 3509 86 3513
rect 89 3509 93 3513
rect 95 3509 99 3513
rect 20 3502 24 3506
rect 38 3502 42 3506
rect 64 3503 68 3507
rect 70 3503 74 3507
rect 76 3503 80 3507
rect 82 3503 86 3507
rect 89 3503 93 3507
rect 95 3503 99 3507
rect 20 3496 24 3500
rect 38 3496 42 3500
rect 64 3497 68 3501
rect 70 3497 74 3501
rect 76 3497 80 3501
rect 82 3497 86 3501
rect 89 3497 93 3501
rect 95 3497 99 3501
rect 20 3490 24 3494
rect 38 3490 42 3494
rect 64 3491 68 3495
rect 70 3491 74 3495
rect 76 3491 80 3495
rect 82 3491 86 3495
rect 89 3491 93 3495
rect 95 3491 99 3495
rect 112 3514 116 3518
rect 125 3514 129 3518
rect 112 3508 116 3512
rect 125 3508 129 3512
rect 112 3502 116 3506
rect 125 3502 129 3506
rect 112 3496 116 3500
rect 125 3496 129 3500
rect 112 3490 116 3494
rect 125 3490 129 3494
rect 20 3142 24 3146
rect 38 3142 42 3146
rect 64 3141 68 3145
rect 70 3141 74 3145
rect 76 3141 80 3145
rect 82 3141 86 3145
rect 89 3141 93 3145
rect 95 3141 99 3145
rect 20 3136 24 3140
rect 38 3136 42 3140
rect 64 3135 68 3139
rect 70 3135 74 3139
rect 76 3135 80 3139
rect 82 3135 86 3139
rect 89 3135 93 3139
rect 95 3135 99 3139
rect 20 3130 24 3134
rect 38 3130 42 3134
rect 64 3129 68 3133
rect 70 3129 74 3133
rect 76 3129 80 3133
rect 82 3129 86 3133
rect 89 3129 93 3133
rect 95 3129 99 3133
rect 20 3124 24 3128
rect 38 3124 42 3128
rect 64 3123 68 3127
rect 70 3123 74 3127
rect 76 3123 80 3127
rect 82 3123 86 3127
rect 89 3123 93 3127
rect 95 3123 99 3127
rect 20 3118 24 3122
rect 38 3118 42 3122
rect 64 3117 68 3121
rect 70 3117 74 3121
rect 76 3117 80 3121
rect 82 3117 86 3121
rect 89 3117 93 3121
rect 95 3117 99 3121
rect 112 3142 116 3146
rect 125 3142 129 3146
rect 112 3136 116 3140
rect 125 3136 129 3140
rect 112 3130 116 3134
rect 125 3130 129 3134
rect 112 3124 116 3128
rect 125 3124 129 3128
rect 112 3118 116 3122
rect 125 3118 129 3122
rect 20 3112 24 3116
rect 38 3112 42 3116
rect 112 3112 116 3116
rect 125 3112 129 3116
rect 20 3106 24 3110
rect 38 3106 42 3110
rect 53 3108 57 3112
rect 112 3106 116 3110
rect 125 3106 129 3110
rect 53 3098 57 3102
rect 53 3060 57 3064
rect 20 3052 24 3056
rect 38 3052 42 3056
rect 53 3050 57 3054
rect 112 3052 116 3056
rect 125 3052 129 3056
rect 20 3046 24 3050
rect 38 3046 42 3050
rect 112 3046 116 3050
rect 125 3046 129 3050
rect 20 3040 24 3044
rect 38 3040 42 3044
rect 64 3041 68 3045
rect 70 3041 74 3045
rect 76 3041 80 3045
rect 82 3041 86 3045
rect 89 3041 93 3045
rect 95 3041 99 3045
rect 20 3034 24 3038
rect 38 3034 42 3038
rect 64 3035 68 3039
rect 70 3035 74 3039
rect 76 3035 80 3039
rect 82 3035 86 3039
rect 89 3035 93 3039
rect 95 3035 99 3039
rect 20 3028 24 3032
rect 38 3028 42 3032
rect 64 3029 68 3033
rect 70 3029 74 3033
rect 76 3029 80 3033
rect 82 3029 86 3033
rect 89 3029 93 3033
rect 95 3029 99 3033
rect 20 3022 24 3026
rect 38 3022 42 3026
rect 64 3023 68 3027
rect 70 3023 74 3027
rect 76 3023 80 3027
rect 82 3023 86 3027
rect 89 3023 93 3027
rect 95 3023 99 3027
rect 20 3016 24 3020
rect 38 3016 42 3020
rect 64 3017 68 3021
rect 70 3017 74 3021
rect 76 3017 80 3021
rect 82 3017 86 3021
rect 89 3017 93 3021
rect 95 3017 99 3021
rect 112 3040 116 3044
rect 125 3040 129 3044
rect 112 3034 116 3038
rect 125 3034 129 3038
rect 112 3028 116 3032
rect 125 3028 129 3032
rect 112 3022 116 3026
rect 125 3022 129 3026
rect 112 3016 116 3020
rect 125 3016 129 3020
rect 20 2668 24 2672
rect 38 2668 42 2672
rect 64 2667 68 2671
rect 70 2667 74 2671
rect 76 2667 80 2671
rect 82 2667 86 2671
rect 89 2667 93 2671
rect 95 2667 99 2671
rect 20 2662 24 2666
rect 38 2662 42 2666
rect 64 2661 68 2665
rect 70 2661 74 2665
rect 76 2661 80 2665
rect 82 2661 86 2665
rect 89 2661 93 2665
rect 95 2661 99 2665
rect 20 2656 24 2660
rect 38 2656 42 2660
rect 64 2655 68 2659
rect 70 2655 74 2659
rect 76 2655 80 2659
rect 82 2655 86 2659
rect 89 2655 93 2659
rect 95 2655 99 2659
rect 20 2650 24 2654
rect 38 2650 42 2654
rect 64 2649 68 2653
rect 70 2649 74 2653
rect 76 2649 80 2653
rect 82 2649 86 2653
rect 89 2649 93 2653
rect 95 2649 99 2653
rect 20 2644 24 2648
rect 38 2644 42 2648
rect 64 2643 68 2647
rect 70 2643 74 2647
rect 76 2643 80 2647
rect 82 2643 86 2647
rect 89 2643 93 2647
rect 95 2643 99 2647
rect 112 2668 116 2672
rect 125 2668 129 2672
rect 112 2662 116 2666
rect 125 2662 129 2666
rect 112 2656 116 2660
rect 125 2656 129 2660
rect 112 2650 116 2654
rect 125 2650 129 2654
rect 112 2644 116 2648
rect 125 2644 129 2648
rect 20 2638 24 2642
rect 38 2638 42 2642
rect 112 2638 116 2642
rect 125 2638 129 2642
rect 20 2632 24 2636
rect 38 2632 42 2636
rect 53 2634 57 2638
rect 112 2632 116 2636
rect 125 2632 129 2636
rect 53 2624 57 2628
rect 53 2586 57 2590
rect 20 2578 24 2582
rect 38 2578 42 2582
rect 53 2576 57 2580
rect 112 2578 116 2582
rect 125 2578 129 2582
rect 20 2572 24 2576
rect 38 2572 42 2576
rect 112 2572 116 2576
rect 125 2572 129 2576
rect 20 2566 24 2570
rect 38 2566 42 2570
rect 64 2567 68 2571
rect 70 2567 74 2571
rect 76 2567 80 2571
rect 82 2567 86 2571
rect 89 2567 93 2571
rect 95 2567 99 2571
rect 20 2560 24 2564
rect 38 2560 42 2564
rect 64 2561 68 2565
rect 70 2561 74 2565
rect 76 2561 80 2565
rect 82 2561 86 2565
rect 89 2561 93 2565
rect 95 2561 99 2565
rect 20 2554 24 2558
rect 38 2554 42 2558
rect 64 2555 68 2559
rect 70 2555 74 2559
rect 76 2555 80 2559
rect 82 2555 86 2559
rect 89 2555 93 2559
rect 95 2555 99 2559
rect 20 2548 24 2552
rect 38 2548 42 2552
rect 64 2549 68 2553
rect 70 2549 74 2553
rect 76 2549 80 2553
rect 82 2549 86 2553
rect 89 2549 93 2553
rect 95 2549 99 2553
rect 20 2542 24 2546
rect 38 2542 42 2546
rect 64 2543 68 2547
rect 70 2543 74 2547
rect 76 2543 80 2547
rect 82 2543 86 2547
rect 89 2543 93 2547
rect 95 2543 99 2547
rect 112 2566 116 2570
rect 125 2566 129 2570
rect 112 2560 116 2564
rect 125 2560 129 2564
rect 112 2554 116 2558
rect 125 2554 129 2558
rect 112 2548 116 2552
rect 125 2548 129 2552
rect 112 2542 116 2546
rect 125 2542 129 2546
rect 20 2194 24 2198
rect 38 2194 42 2198
rect 64 2193 68 2197
rect 70 2193 74 2197
rect 76 2193 80 2197
rect 82 2193 86 2197
rect 89 2193 93 2197
rect 95 2193 99 2197
rect 20 2188 24 2192
rect 38 2188 42 2192
rect 64 2187 68 2191
rect 70 2187 74 2191
rect 76 2187 80 2191
rect 82 2187 86 2191
rect 89 2187 93 2191
rect 95 2187 99 2191
rect 20 2182 24 2186
rect 38 2182 42 2186
rect 64 2181 68 2185
rect 70 2181 74 2185
rect 76 2181 80 2185
rect 82 2181 86 2185
rect 89 2181 93 2185
rect 95 2181 99 2185
rect 20 2176 24 2180
rect 38 2176 42 2180
rect 64 2175 68 2179
rect 70 2175 74 2179
rect 76 2175 80 2179
rect 82 2175 86 2179
rect 89 2175 93 2179
rect 95 2175 99 2179
rect 20 2170 24 2174
rect 38 2170 42 2174
rect 64 2169 68 2173
rect 70 2169 74 2173
rect 76 2169 80 2173
rect 82 2169 86 2173
rect 89 2169 93 2173
rect 95 2169 99 2173
rect 112 2194 116 2198
rect 125 2194 129 2198
rect 112 2188 116 2192
rect 125 2188 129 2192
rect 112 2182 116 2186
rect 125 2182 129 2186
rect 112 2176 116 2180
rect 125 2176 129 2180
rect 112 2170 116 2174
rect 125 2170 129 2174
rect 20 2164 24 2168
rect 38 2164 42 2168
rect 112 2164 116 2168
rect 125 2164 129 2168
rect 20 2158 24 2162
rect 38 2158 42 2162
rect 53 2160 57 2164
rect 112 2158 116 2162
rect 125 2158 129 2162
rect 53 2150 57 2154
rect 53 2112 57 2116
rect 20 2104 24 2108
rect 38 2104 42 2108
rect 53 2102 57 2106
rect 112 2104 116 2108
rect 125 2104 129 2108
rect 20 2098 24 2102
rect 38 2098 42 2102
rect 112 2098 116 2102
rect 125 2098 129 2102
rect 20 2092 24 2096
rect 38 2092 42 2096
rect 64 2093 68 2097
rect 70 2093 74 2097
rect 76 2093 80 2097
rect 82 2093 86 2097
rect 89 2093 93 2097
rect 95 2093 99 2097
rect 20 2086 24 2090
rect 38 2086 42 2090
rect 64 2087 68 2091
rect 70 2087 74 2091
rect 76 2087 80 2091
rect 82 2087 86 2091
rect 89 2087 93 2091
rect 95 2087 99 2091
rect 20 2080 24 2084
rect 38 2080 42 2084
rect 64 2081 68 2085
rect 70 2081 74 2085
rect 76 2081 80 2085
rect 82 2081 86 2085
rect 89 2081 93 2085
rect 95 2081 99 2085
rect 20 2074 24 2078
rect 38 2074 42 2078
rect 64 2075 68 2079
rect 70 2075 74 2079
rect 76 2075 80 2079
rect 82 2075 86 2079
rect 89 2075 93 2079
rect 95 2075 99 2079
rect 20 2068 24 2072
rect 38 2068 42 2072
rect 64 2069 68 2073
rect 70 2069 74 2073
rect 76 2069 80 2073
rect 82 2069 86 2073
rect 89 2069 93 2073
rect 95 2069 99 2073
rect 112 2092 116 2096
rect 125 2092 129 2096
rect 112 2086 116 2090
rect 125 2086 129 2090
rect 112 2080 116 2084
rect 125 2080 129 2084
rect 112 2074 116 2078
rect 125 2074 129 2078
rect 112 2068 116 2072
rect 125 2068 129 2072
rect 20 1720 24 1724
rect 38 1720 42 1724
rect 64 1719 68 1723
rect 70 1719 74 1723
rect 76 1719 80 1723
rect 82 1719 86 1723
rect 89 1719 93 1723
rect 95 1719 99 1723
rect 20 1714 24 1718
rect 38 1714 42 1718
rect 64 1713 68 1717
rect 70 1713 74 1717
rect 76 1713 80 1717
rect 82 1713 86 1717
rect 89 1713 93 1717
rect 95 1713 99 1717
rect 20 1708 24 1712
rect 38 1708 42 1712
rect 64 1707 68 1711
rect 70 1707 74 1711
rect 76 1707 80 1711
rect 82 1707 86 1711
rect 89 1707 93 1711
rect 95 1707 99 1711
rect 20 1702 24 1706
rect 38 1702 42 1706
rect 64 1701 68 1705
rect 70 1701 74 1705
rect 76 1701 80 1705
rect 82 1701 86 1705
rect 89 1701 93 1705
rect 95 1701 99 1705
rect 20 1696 24 1700
rect 38 1696 42 1700
rect 64 1695 68 1699
rect 70 1695 74 1699
rect 76 1695 80 1699
rect 82 1695 86 1699
rect 89 1695 93 1699
rect 95 1695 99 1699
rect 112 1720 116 1724
rect 125 1720 129 1724
rect 112 1714 116 1718
rect 125 1714 129 1718
rect 112 1708 116 1712
rect 125 1708 129 1712
rect 112 1702 116 1706
rect 125 1702 129 1706
rect 112 1696 116 1700
rect 125 1696 129 1700
rect 20 1690 24 1694
rect 38 1690 42 1694
rect 112 1690 116 1694
rect 125 1690 129 1694
rect 20 1684 24 1688
rect 38 1684 42 1688
rect 53 1686 57 1690
rect 112 1684 116 1688
rect 125 1684 129 1688
rect 53 1676 57 1680
rect 53 1638 57 1642
rect 20 1630 24 1634
rect 38 1630 42 1634
rect 53 1628 57 1632
rect 112 1630 116 1634
rect 125 1630 129 1634
rect 20 1624 24 1628
rect 38 1624 42 1628
rect 112 1624 116 1628
rect 125 1624 129 1628
rect 20 1618 24 1622
rect 38 1618 42 1622
rect 64 1619 68 1623
rect 70 1619 74 1623
rect 76 1619 80 1623
rect 82 1619 86 1623
rect 89 1619 93 1623
rect 95 1619 99 1623
rect 20 1612 24 1616
rect 38 1612 42 1616
rect 64 1613 68 1617
rect 70 1613 74 1617
rect 76 1613 80 1617
rect 82 1613 86 1617
rect 89 1613 93 1617
rect 95 1613 99 1617
rect 20 1606 24 1610
rect 38 1606 42 1610
rect 64 1607 68 1611
rect 70 1607 74 1611
rect 76 1607 80 1611
rect 82 1607 86 1611
rect 89 1607 93 1611
rect 95 1607 99 1611
rect 20 1600 24 1604
rect 38 1600 42 1604
rect 64 1601 68 1605
rect 70 1601 74 1605
rect 76 1601 80 1605
rect 82 1601 86 1605
rect 89 1601 93 1605
rect 95 1601 99 1605
rect 20 1594 24 1598
rect 38 1594 42 1598
rect 64 1595 68 1599
rect 70 1595 74 1599
rect 76 1595 80 1599
rect 82 1595 86 1599
rect 89 1595 93 1599
rect 95 1595 99 1599
rect 112 1618 116 1622
rect 125 1618 129 1622
rect 112 1612 116 1616
rect 125 1612 129 1616
rect 112 1606 116 1610
rect 125 1606 129 1610
rect 112 1600 116 1604
rect 125 1600 129 1604
rect 112 1594 116 1598
rect 125 1594 129 1598
rect 20 1246 24 1250
rect 38 1246 42 1250
rect 64 1245 68 1249
rect 70 1245 74 1249
rect 76 1245 80 1249
rect 82 1245 86 1249
rect 89 1245 93 1249
rect 95 1245 99 1249
rect 20 1240 24 1244
rect 38 1240 42 1244
rect 64 1239 68 1243
rect 70 1239 74 1243
rect 76 1239 80 1243
rect 82 1239 86 1243
rect 89 1239 93 1243
rect 95 1239 99 1243
rect 20 1234 24 1238
rect 38 1234 42 1238
rect 64 1233 68 1237
rect 70 1233 74 1237
rect 76 1233 80 1237
rect 82 1233 86 1237
rect 89 1233 93 1237
rect 95 1233 99 1237
rect 20 1228 24 1232
rect 38 1228 42 1232
rect 64 1227 68 1231
rect 70 1227 74 1231
rect 76 1227 80 1231
rect 82 1227 86 1231
rect 89 1227 93 1231
rect 95 1227 99 1231
rect 20 1222 24 1226
rect 38 1222 42 1226
rect 64 1221 68 1225
rect 70 1221 74 1225
rect 76 1221 80 1225
rect 82 1221 86 1225
rect 89 1221 93 1225
rect 95 1221 99 1225
rect 112 1246 116 1250
rect 125 1246 129 1250
rect 112 1240 116 1244
rect 125 1240 129 1244
rect 112 1234 116 1238
rect 125 1234 129 1238
rect 112 1228 116 1232
rect 125 1228 129 1232
rect 112 1222 116 1226
rect 125 1222 129 1226
rect 20 1216 24 1220
rect 38 1216 42 1220
rect 112 1216 116 1220
rect 125 1216 129 1220
rect 20 1210 24 1214
rect 38 1210 42 1214
rect 53 1212 57 1216
rect 112 1210 116 1214
rect 125 1210 129 1214
rect 53 1202 57 1206
rect 53 1164 57 1168
rect 20 1156 24 1160
rect 38 1156 42 1160
rect 53 1154 57 1158
rect 112 1156 116 1160
rect 125 1156 129 1160
rect 20 1150 24 1154
rect 38 1150 42 1154
rect 112 1150 116 1154
rect 125 1150 129 1154
rect 20 1144 24 1148
rect 38 1144 42 1148
rect 64 1145 68 1149
rect 70 1145 74 1149
rect 76 1145 80 1149
rect 82 1145 86 1149
rect 89 1145 93 1149
rect 95 1145 99 1149
rect 20 1138 24 1142
rect 38 1138 42 1142
rect 64 1139 68 1143
rect 70 1139 74 1143
rect 76 1139 80 1143
rect 82 1139 86 1143
rect 89 1139 93 1143
rect 95 1139 99 1143
rect 20 1132 24 1136
rect 38 1132 42 1136
rect 64 1133 68 1137
rect 70 1133 74 1137
rect 76 1133 80 1137
rect 82 1133 86 1137
rect 89 1133 93 1137
rect 95 1133 99 1137
rect 20 1126 24 1130
rect 38 1126 42 1130
rect 64 1127 68 1131
rect 70 1127 74 1131
rect 76 1127 80 1131
rect 82 1127 86 1131
rect 89 1127 93 1131
rect 95 1127 99 1131
rect 20 1120 24 1124
rect 38 1120 42 1124
rect 64 1121 68 1125
rect 70 1121 74 1125
rect 76 1121 80 1125
rect 82 1121 86 1125
rect 89 1121 93 1125
rect 95 1121 99 1125
rect 112 1144 116 1148
rect 125 1144 129 1148
rect 112 1138 116 1142
rect 125 1138 129 1142
rect 112 1132 116 1136
rect 125 1132 129 1136
rect 112 1126 116 1130
rect 125 1126 129 1130
rect 112 1120 116 1124
rect 125 1120 129 1124
rect 20 772 24 776
rect 38 772 42 776
rect 64 771 68 775
rect 70 771 74 775
rect 76 771 80 775
rect 82 771 86 775
rect 89 771 93 775
rect 95 771 99 775
rect 20 766 24 770
rect 38 766 42 770
rect 64 765 68 769
rect 70 765 74 769
rect 76 765 80 769
rect 82 765 86 769
rect 89 765 93 769
rect 95 765 99 769
rect 20 760 24 764
rect 38 760 42 764
rect 64 759 68 763
rect 70 759 74 763
rect 76 759 80 763
rect 82 759 86 763
rect 89 759 93 763
rect 95 759 99 763
rect 20 754 24 758
rect 38 754 42 758
rect 64 753 68 757
rect 70 753 74 757
rect 76 753 80 757
rect 82 753 86 757
rect 89 753 93 757
rect 95 753 99 757
rect 20 748 24 752
rect 38 748 42 752
rect 64 747 68 751
rect 70 747 74 751
rect 76 747 80 751
rect 82 747 86 751
rect 89 747 93 751
rect 95 747 99 751
rect 112 772 116 776
rect 125 772 129 776
rect 112 766 116 770
rect 125 766 129 770
rect 112 760 116 764
rect 125 760 129 764
rect 112 754 116 758
rect 125 754 129 758
rect 112 748 116 752
rect 125 748 129 752
rect 20 742 24 746
rect 38 742 42 746
rect 112 742 116 746
rect 125 742 129 746
rect 20 736 24 740
rect 38 736 42 740
rect 53 738 57 742
rect 112 736 116 740
rect 125 736 129 740
rect 53 728 57 732
rect 53 690 57 694
rect 20 682 24 686
rect 38 682 42 686
rect 53 680 57 684
rect 112 682 116 686
rect 125 682 129 686
rect 20 676 24 680
rect 38 676 42 680
rect 112 676 116 680
rect 125 676 129 680
rect 20 670 24 674
rect 38 670 42 674
rect 64 671 68 675
rect 70 671 74 675
rect 76 671 80 675
rect 82 671 86 675
rect 89 671 93 675
rect 95 671 99 675
rect 20 664 24 668
rect 38 664 42 668
rect 64 665 68 669
rect 70 665 74 669
rect 76 665 80 669
rect 82 665 86 669
rect 89 665 93 669
rect 95 665 99 669
rect 20 658 24 662
rect 38 658 42 662
rect 64 659 68 663
rect 70 659 74 663
rect 76 659 80 663
rect 82 659 86 663
rect 89 659 93 663
rect 95 659 99 663
rect 20 652 24 656
rect 38 652 42 656
rect 64 653 68 657
rect 70 653 74 657
rect 76 653 80 657
rect 82 653 86 657
rect 89 653 93 657
rect 95 653 99 657
rect 20 646 24 650
rect 38 646 42 650
rect 64 647 68 651
rect 70 647 74 651
rect 76 647 80 651
rect 82 647 86 651
rect 89 647 93 651
rect 95 647 99 651
rect 112 670 116 674
rect 125 670 129 674
rect 112 664 116 668
rect 125 664 129 668
rect 112 658 116 662
rect 125 658 129 662
rect 112 652 116 656
rect 125 652 129 656
rect 112 646 116 650
rect 125 646 129 650
rect 20 298 24 302
rect 38 298 42 302
rect 64 297 68 301
rect 70 297 74 301
rect 76 297 80 301
rect 82 297 86 301
rect 89 297 93 301
rect 95 297 99 301
rect 20 292 24 296
rect 38 292 42 296
rect 64 291 68 295
rect 70 291 74 295
rect 76 291 80 295
rect 82 291 86 295
rect 89 291 93 295
rect 95 291 99 295
rect 20 286 24 290
rect 38 286 42 290
rect 64 285 68 289
rect 70 285 74 289
rect 76 285 80 289
rect 82 285 86 289
rect 89 285 93 289
rect 95 285 99 289
rect 20 280 24 284
rect 38 280 42 284
rect 64 279 68 283
rect 70 279 74 283
rect 76 279 80 283
rect 82 279 86 283
rect 89 279 93 283
rect 95 279 99 283
rect 20 274 24 278
rect 38 274 42 278
rect 64 273 68 277
rect 70 273 74 277
rect 76 273 80 277
rect 82 273 86 277
rect 89 273 93 277
rect 95 273 99 277
rect 112 298 116 302
rect 125 298 129 302
rect 112 292 116 296
rect 125 292 129 296
rect 112 286 116 290
rect 125 286 129 290
rect 112 280 116 284
rect 125 280 129 284
rect 112 274 116 278
rect 125 274 129 278
rect 20 268 24 272
rect 38 268 42 272
rect 112 268 116 272
rect 125 268 129 272
rect 20 262 24 266
rect 38 262 42 266
rect 53 264 57 268
rect 112 262 116 266
rect 125 262 129 266
rect 53 254 57 258
rect 53 216 57 220
rect 20 208 24 212
rect 38 208 42 212
rect 53 206 57 210
rect 112 208 116 212
rect 125 208 129 212
rect 20 202 24 206
rect 38 202 42 206
rect 112 202 116 206
rect 125 202 129 206
rect 20 196 24 200
rect 38 196 42 200
rect 64 197 68 201
rect 70 197 74 201
rect 76 197 80 201
rect 82 197 86 201
rect 89 197 93 201
rect 95 197 99 201
rect 20 190 24 194
rect 38 190 42 194
rect 64 191 68 195
rect 70 191 74 195
rect 76 191 80 195
rect 82 191 86 195
rect 89 191 93 195
rect 95 191 99 195
rect 20 184 24 188
rect 38 184 42 188
rect 64 185 68 189
rect 70 185 74 189
rect 76 185 80 189
rect 82 185 86 189
rect 89 185 93 189
rect 95 185 99 189
rect 20 178 24 182
rect 38 178 42 182
rect 64 179 68 183
rect 70 179 74 183
rect 76 179 80 183
rect 82 179 86 183
rect 89 179 93 183
rect 95 179 99 183
rect 20 172 24 176
rect 38 172 42 176
rect 64 173 68 177
rect 70 173 74 177
rect 76 173 80 177
rect 82 173 86 177
rect 89 173 93 177
rect 95 173 99 177
rect 112 196 116 200
rect 125 196 129 200
rect 112 190 116 194
rect 125 190 129 194
rect 112 184 116 188
rect 125 184 129 188
rect 112 178 116 182
rect 125 178 129 182
rect 112 172 116 176
rect 125 172 129 176
<< electrodecap >>
rect 12 3965 48 4168
rect 17 3915 48 3965
rect 12 3669 48 3915
rect 17 3619 48 3669
rect 12 3491 48 3619
rect 17 3441 48 3491
rect 12 3195 48 3441
rect 17 3145 48 3195
rect 12 3017 48 3145
rect 17 2967 48 3017
rect 12 2721 48 2967
rect 17 2671 48 2721
rect 12 2543 48 2671
rect 17 2493 48 2543
rect 12 2247 48 2493
rect 17 2197 48 2247
rect 12 2069 48 2197
rect 17 2019 48 2069
rect 12 1773 48 2019
rect 17 1723 48 1773
rect 12 1595 48 1723
rect 17 1545 48 1595
rect 12 1299 48 1545
rect 17 1249 48 1299
rect 12 1121 48 1249
rect 17 1071 48 1121
rect 12 825 48 1071
rect 17 775 48 825
rect 12 647 48 775
rect 17 597 48 647
rect 12 351 48 597
rect 17 301 48 351
rect 12 98 48 301
rect 51 95 59 4171
rect 62 84 102 4182
rect 105 4143 137 4257
rect 105 4093 132 4143
rect 105 3965 137 4093
rect 105 3915 132 3965
rect 105 3669 137 3915
rect 105 3619 132 3669
rect 105 3491 137 3619
rect 105 3441 132 3491
rect 105 3195 137 3441
rect 105 3145 132 3195
rect 105 3017 137 3145
rect 105 2967 132 3017
rect 105 2721 137 2967
rect 105 2671 132 2721
rect 105 2543 137 2671
rect 105 2493 132 2543
rect 105 2247 137 2493
rect 105 2197 132 2247
rect 105 2069 137 2197
rect 105 2019 132 2069
rect 105 1773 137 2019
rect 105 1723 132 1773
rect 105 1595 137 1723
rect 105 1545 132 1595
rect 105 1299 137 1545
rect 105 1249 132 1299
rect 105 1121 137 1249
rect 105 1071 132 1121
rect 105 825 137 1071
rect 105 775 132 825
rect 105 647 137 775
rect 105 597 132 647
rect 105 351 137 597
rect 105 301 132 351
rect 105 173 137 301
rect 105 123 132 173
rect 105 41 137 123
<< psubstratepdiff >>
rect 143 4262 149 4263
rect 143 4258 144 4262
rect 148 4258 149 4262
rect 143 4256 149 4258
rect 143 4252 144 4256
rect 148 4252 149 4256
rect 143 4250 149 4252
rect 143 4246 144 4250
rect 148 4246 149 4250
rect 143 4244 149 4246
rect 143 4240 144 4244
rect 148 4240 149 4244
rect 143 4238 149 4240
rect 143 4234 144 4238
rect 148 4234 149 4238
rect 143 4232 149 4234
rect 143 4228 144 4232
rect 148 4228 149 4232
rect 143 4226 149 4228
rect 143 4222 144 4226
rect 148 4222 149 4226
rect 143 4220 149 4222
rect 143 4216 144 4220
rect 148 4216 149 4220
rect 143 4214 149 4216
rect 143 4210 144 4214
rect 148 4210 149 4214
rect 143 4208 149 4210
rect 143 4204 144 4208
rect 148 4204 149 4208
rect 143 4202 149 4204
rect 143 4198 144 4202
rect 148 4198 149 4202
rect 143 4196 149 4198
rect 143 4192 144 4196
rect 148 4192 149 4196
rect 143 4190 149 4192
rect 143 4186 144 4190
rect 148 4186 149 4190
rect 143 4184 149 4186
rect 143 4180 144 4184
rect 148 4180 149 4184
rect 143 4178 149 4180
rect 143 4174 144 4178
rect 148 4174 149 4178
rect 143 4172 149 4174
rect 143 4168 144 4172
rect 148 4168 149 4172
rect 143 4166 149 4168
rect 143 4162 144 4166
rect 148 4162 149 4166
rect 143 4160 149 4162
rect 143 4156 144 4160
rect 148 4156 149 4160
rect 143 4154 149 4156
rect 143 4150 144 4154
rect 148 4150 149 4154
rect 143 4148 149 4150
rect 143 4144 144 4148
rect 148 4144 149 4148
rect 143 4142 149 4144
rect 143 4138 144 4142
rect 148 4138 149 4142
rect 143 4136 149 4138
rect 143 4132 144 4136
rect 148 4132 149 4136
rect 143 4130 149 4132
rect 143 4126 144 4130
rect 148 4126 149 4130
rect 143 4124 149 4126
rect 143 4120 144 4124
rect 148 4120 149 4124
rect 143 4118 149 4120
rect 143 4114 144 4118
rect 148 4114 149 4118
rect 143 4112 149 4114
rect 143 4108 144 4112
rect 148 4108 149 4112
rect 143 4106 149 4108
rect 143 4102 144 4106
rect 148 4102 149 4106
rect 143 4100 149 4102
rect 143 4096 144 4100
rect 148 4096 149 4100
rect 143 4094 149 4096
rect 143 4090 144 4094
rect 148 4090 149 4094
rect 143 4088 149 4090
rect 143 4084 144 4088
rect 148 4084 149 4088
rect 143 4082 149 4084
rect 143 4078 144 4082
rect 148 4078 149 4082
rect 143 4076 149 4078
rect 143 4072 144 4076
rect 148 4072 149 4076
rect 143 4070 149 4072
rect 143 4066 144 4070
rect 148 4066 149 4070
rect 143 4064 149 4066
rect 143 4060 144 4064
rect 148 4060 149 4064
rect 143 4058 149 4060
rect 143 4054 144 4058
rect 148 4054 149 4058
rect 143 4052 149 4054
rect 143 4048 144 4052
rect 148 4048 149 4052
rect 143 4046 149 4048
rect 143 4042 144 4046
rect 148 4042 149 4046
rect 143 4016 149 4042
rect 143 4012 144 4016
rect 148 4012 149 4016
rect 143 4010 149 4012
rect 143 4006 144 4010
rect 148 4006 149 4010
rect 143 4004 149 4006
rect 143 4000 144 4004
rect 148 4000 149 4004
rect 143 3998 149 4000
rect 143 3994 144 3998
rect 148 3994 149 3998
rect 143 3992 149 3994
rect 143 3988 144 3992
rect 148 3988 149 3992
rect 143 3986 149 3988
rect 143 3982 144 3986
rect 148 3982 149 3986
rect 143 3980 149 3982
rect 143 3976 144 3980
rect 148 3976 149 3980
rect 143 3974 149 3976
rect 143 3970 144 3974
rect 148 3970 149 3974
rect 143 3968 149 3970
rect 143 3964 144 3968
rect 148 3964 149 3968
rect 143 3962 149 3964
rect 143 3958 144 3962
rect 148 3958 149 3962
rect 143 3956 149 3958
rect 143 3952 144 3956
rect 148 3952 149 3956
rect 143 3950 149 3952
rect 143 3946 144 3950
rect 148 3946 149 3950
rect 143 3944 149 3946
rect 143 3940 144 3944
rect 148 3940 149 3944
rect 143 3938 149 3940
rect 143 3934 144 3938
rect 148 3934 149 3938
rect 143 3932 149 3934
rect 143 3928 144 3932
rect 148 3928 149 3932
rect 143 3926 149 3928
rect 143 3922 144 3926
rect 148 3922 149 3926
rect 143 3920 149 3922
rect 143 3916 144 3920
rect 148 3916 149 3920
rect 143 3914 149 3916
rect 143 3910 144 3914
rect 148 3910 149 3914
rect 143 3908 149 3910
rect 143 3904 144 3908
rect 148 3904 149 3908
rect 143 3902 149 3904
rect 143 3898 144 3902
rect 148 3898 149 3902
rect 143 3896 149 3898
rect 143 3892 144 3896
rect 148 3892 149 3896
rect 143 3890 149 3892
rect 143 3886 144 3890
rect 148 3886 149 3890
rect 143 3884 149 3886
rect 143 3880 144 3884
rect 148 3880 149 3884
rect 143 3878 149 3880
rect 143 3874 144 3878
rect 148 3874 149 3878
rect 143 3872 149 3874
rect 143 3868 144 3872
rect 148 3868 149 3872
rect 143 3866 149 3868
rect 143 3862 144 3866
rect 148 3862 149 3866
rect 143 3860 149 3862
rect 143 3856 144 3860
rect 148 3856 149 3860
rect 143 3854 149 3856
rect 143 3850 144 3854
rect 148 3850 149 3854
rect 143 3848 149 3850
rect 143 3844 144 3848
rect 148 3844 149 3848
rect 143 3842 149 3844
rect 143 3838 144 3842
rect 148 3838 149 3842
rect 143 3836 149 3838
rect 143 3832 144 3836
rect 148 3832 149 3836
rect 143 3830 149 3832
rect 143 3826 144 3830
rect 148 3826 149 3830
rect 143 3824 149 3826
rect 143 3820 144 3824
rect 148 3820 149 3824
rect 143 3818 149 3820
rect 143 3814 144 3818
rect 148 3814 149 3818
rect 143 3812 149 3814
rect 143 3808 144 3812
rect 148 3808 149 3812
rect 143 3806 149 3808
rect 143 3802 144 3806
rect 148 3802 149 3806
rect 143 3800 149 3802
rect 143 3796 144 3800
rect 148 3796 149 3800
rect 143 3795 149 3796
rect 143 3794 511 3795
rect 143 3790 144 3794
rect 148 3790 150 3794
rect 154 3790 156 3794
rect 160 3790 162 3794
rect 166 3790 168 3794
rect 172 3790 174 3794
rect 178 3790 180 3794
rect 184 3790 186 3794
rect 190 3790 192 3794
rect 196 3790 198 3794
rect 202 3790 204 3794
rect 208 3790 210 3794
rect 214 3790 216 3794
rect 220 3790 222 3794
rect 226 3790 228 3794
rect 232 3790 234 3794
rect 238 3790 240 3794
rect 244 3790 246 3794
rect 250 3790 252 3794
rect 256 3790 258 3794
rect 262 3790 264 3794
rect 268 3790 270 3794
rect 274 3790 276 3794
rect 280 3790 282 3794
rect 286 3790 288 3794
rect 292 3790 294 3794
rect 298 3790 300 3794
rect 304 3790 306 3794
rect 310 3790 312 3794
rect 316 3790 318 3794
rect 322 3790 324 3794
rect 328 3790 330 3794
rect 334 3790 336 3794
rect 340 3790 342 3794
rect 346 3790 348 3794
rect 352 3790 354 3794
rect 358 3790 360 3794
rect 364 3790 366 3794
rect 370 3790 372 3794
rect 376 3790 378 3794
rect 382 3790 384 3794
rect 388 3790 390 3794
rect 394 3790 396 3794
rect 400 3790 402 3794
rect 406 3790 408 3794
rect 412 3790 414 3794
rect 418 3790 420 3794
rect 424 3790 426 3794
rect 430 3790 432 3794
rect 436 3790 438 3794
rect 442 3790 444 3794
rect 448 3790 450 3794
rect 454 3790 456 3794
rect 460 3790 462 3794
rect 466 3790 468 3794
rect 472 3790 474 3794
rect 478 3790 480 3794
rect 484 3790 486 3794
rect 490 3790 492 3794
rect 496 3790 498 3794
rect 502 3790 504 3794
rect 508 3790 511 3794
rect 143 3789 511 3790
rect 143 3788 149 3789
rect 143 3784 144 3788
rect 148 3784 149 3788
rect 143 3782 149 3784
rect 143 3778 144 3782
rect 148 3778 149 3782
rect 143 3776 149 3778
rect 143 3772 144 3776
rect 148 3772 149 3776
rect 143 3770 149 3772
rect 143 3766 144 3770
rect 148 3766 149 3770
rect 143 3764 149 3766
rect 143 3760 144 3764
rect 148 3760 149 3764
rect 143 3758 149 3760
rect 143 3754 144 3758
rect 148 3754 149 3758
rect 143 3752 149 3754
rect 143 3748 144 3752
rect 148 3748 149 3752
rect 143 3746 149 3748
rect 143 3742 144 3746
rect 148 3742 149 3746
rect 143 3740 149 3742
rect 143 3736 144 3740
rect 148 3736 149 3740
rect 143 3734 149 3736
rect 143 3730 144 3734
rect 148 3730 149 3734
rect 143 3728 149 3730
rect 143 3724 144 3728
rect 148 3724 149 3728
rect 143 3722 149 3724
rect 143 3718 144 3722
rect 148 3718 149 3722
rect 143 3716 149 3718
rect 143 3712 144 3716
rect 148 3712 149 3716
rect 143 3710 149 3712
rect 143 3706 144 3710
rect 148 3706 149 3710
rect 143 3704 149 3706
rect 143 3700 144 3704
rect 148 3700 149 3704
rect 143 3698 149 3700
rect 143 3694 144 3698
rect 148 3694 149 3698
rect 143 3692 149 3694
rect 143 3688 144 3692
rect 148 3688 149 3692
rect 143 3686 149 3688
rect 143 3682 144 3686
rect 148 3682 149 3686
rect 143 3680 149 3682
rect 143 3676 144 3680
rect 148 3676 149 3680
rect 143 3674 149 3676
rect 143 3670 144 3674
rect 148 3670 149 3674
rect 143 3668 149 3670
rect 143 3664 144 3668
rect 148 3664 149 3668
rect 143 3662 149 3664
rect 143 3658 144 3662
rect 148 3658 149 3662
rect 143 3656 149 3658
rect 143 3652 144 3656
rect 148 3652 149 3656
rect 143 3650 149 3652
rect 143 3646 144 3650
rect 148 3646 149 3650
rect 143 3644 149 3646
rect 143 3640 144 3644
rect 148 3640 149 3644
rect 143 3638 149 3640
rect 143 3634 144 3638
rect 148 3634 149 3638
rect 143 3632 149 3634
rect 143 3628 144 3632
rect 148 3628 149 3632
rect 143 3626 149 3628
rect 143 3622 144 3626
rect 148 3622 149 3626
rect 143 3620 149 3622
rect 143 3616 144 3620
rect 148 3616 149 3620
rect 143 3614 149 3616
rect 143 3610 144 3614
rect 148 3610 149 3614
rect 143 3608 149 3610
rect 143 3604 144 3608
rect 148 3604 149 3608
rect 143 3602 149 3604
rect 143 3598 144 3602
rect 148 3598 149 3602
rect 143 3596 149 3598
rect 143 3592 144 3596
rect 148 3592 149 3596
rect 143 3590 149 3592
rect 143 3586 144 3590
rect 148 3586 149 3590
rect 143 3584 149 3586
rect 143 3580 144 3584
rect 148 3580 149 3584
rect 143 3578 149 3580
rect 143 3574 144 3578
rect 148 3574 149 3578
rect 143 3572 149 3574
rect 143 3568 144 3572
rect 148 3568 149 3572
rect 143 3542 149 3568
rect 143 3538 144 3542
rect 148 3538 149 3542
rect 143 3536 149 3538
rect 143 3532 144 3536
rect 148 3532 149 3536
rect 143 3530 149 3532
rect 143 3526 144 3530
rect 148 3526 149 3530
rect 143 3524 149 3526
rect 143 3520 144 3524
rect 148 3520 149 3524
rect 143 3518 149 3520
rect 143 3514 144 3518
rect 148 3514 149 3518
rect 143 3512 149 3514
rect 143 3508 144 3512
rect 148 3508 149 3512
rect 143 3506 149 3508
rect 143 3502 144 3506
rect 148 3502 149 3506
rect 143 3500 149 3502
rect 143 3496 144 3500
rect 148 3496 149 3500
rect 143 3494 149 3496
rect 143 3490 144 3494
rect 148 3490 149 3494
rect 143 3488 149 3490
rect 143 3484 144 3488
rect 148 3484 149 3488
rect 143 3482 149 3484
rect 143 3478 144 3482
rect 148 3478 149 3482
rect 143 3476 149 3478
rect 143 3472 144 3476
rect 148 3472 149 3476
rect 143 3470 149 3472
rect 143 3466 144 3470
rect 148 3466 149 3470
rect 143 3464 149 3466
rect 143 3460 144 3464
rect 148 3460 149 3464
rect 143 3458 149 3460
rect 143 3454 144 3458
rect 148 3454 149 3458
rect 143 3452 149 3454
rect 143 3448 144 3452
rect 148 3448 149 3452
rect 143 3446 149 3448
rect 143 3442 144 3446
rect 148 3442 149 3446
rect 143 3440 149 3442
rect 143 3436 144 3440
rect 148 3436 149 3440
rect 143 3434 149 3436
rect 143 3430 144 3434
rect 148 3430 149 3434
rect 143 3428 149 3430
rect 143 3424 144 3428
rect 148 3424 149 3428
rect 143 3422 149 3424
rect 143 3418 144 3422
rect 148 3418 149 3422
rect 143 3416 149 3418
rect 143 3412 144 3416
rect 148 3412 149 3416
rect 143 3410 149 3412
rect 143 3406 144 3410
rect 148 3406 149 3410
rect 143 3404 149 3406
rect 143 3400 144 3404
rect 148 3400 149 3404
rect 143 3398 149 3400
rect 143 3394 144 3398
rect 148 3394 149 3398
rect 143 3392 149 3394
rect 143 3388 144 3392
rect 148 3388 149 3392
rect 143 3386 149 3388
rect 143 3382 144 3386
rect 148 3382 149 3386
rect 143 3380 149 3382
rect 143 3376 144 3380
rect 148 3376 149 3380
rect 143 3374 149 3376
rect 143 3370 144 3374
rect 148 3370 149 3374
rect 143 3368 149 3370
rect 143 3364 144 3368
rect 148 3364 149 3368
rect 143 3362 149 3364
rect 143 3358 144 3362
rect 148 3358 149 3362
rect 143 3356 149 3358
rect 143 3352 144 3356
rect 148 3352 149 3356
rect 143 3350 149 3352
rect 143 3346 144 3350
rect 148 3346 149 3350
rect 143 3344 149 3346
rect 143 3340 144 3344
rect 148 3340 149 3344
rect 143 3338 149 3340
rect 143 3334 144 3338
rect 148 3334 149 3338
rect 143 3332 149 3334
rect 143 3328 144 3332
rect 148 3328 149 3332
rect 143 3326 149 3328
rect 143 3322 144 3326
rect 148 3322 149 3326
rect 143 3321 149 3322
rect 143 3320 511 3321
rect 143 3316 144 3320
rect 148 3316 150 3320
rect 154 3316 156 3320
rect 160 3316 162 3320
rect 166 3316 168 3320
rect 172 3316 174 3320
rect 178 3316 180 3320
rect 184 3316 186 3320
rect 190 3316 192 3320
rect 196 3316 198 3320
rect 202 3316 204 3320
rect 208 3316 210 3320
rect 214 3316 216 3320
rect 220 3316 222 3320
rect 226 3316 228 3320
rect 232 3316 234 3320
rect 238 3316 240 3320
rect 244 3316 246 3320
rect 250 3316 252 3320
rect 256 3316 258 3320
rect 262 3316 264 3320
rect 268 3316 270 3320
rect 274 3316 276 3320
rect 280 3316 282 3320
rect 286 3316 288 3320
rect 292 3316 294 3320
rect 298 3316 300 3320
rect 304 3316 306 3320
rect 310 3316 312 3320
rect 316 3316 318 3320
rect 322 3316 324 3320
rect 328 3316 330 3320
rect 334 3316 336 3320
rect 340 3316 342 3320
rect 346 3316 348 3320
rect 352 3316 354 3320
rect 358 3316 360 3320
rect 364 3316 366 3320
rect 370 3316 372 3320
rect 376 3316 378 3320
rect 382 3316 384 3320
rect 388 3316 390 3320
rect 394 3316 396 3320
rect 400 3316 402 3320
rect 406 3316 408 3320
rect 412 3316 414 3320
rect 418 3316 420 3320
rect 424 3316 426 3320
rect 430 3316 432 3320
rect 436 3316 438 3320
rect 442 3316 444 3320
rect 448 3316 450 3320
rect 454 3316 456 3320
rect 460 3316 462 3320
rect 466 3316 468 3320
rect 472 3316 474 3320
rect 478 3316 480 3320
rect 484 3316 486 3320
rect 490 3316 492 3320
rect 496 3316 498 3320
rect 502 3316 504 3320
rect 508 3316 511 3320
rect 143 3315 511 3316
rect 143 3314 149 3315
rect 143 3310 144 3314
rect 148 3310 149 3314
rect 143 3308 149 3310
rect 143 3304 144 3308
rect 148 3304 149 3308
rect 143 3302 149 3304
rect 143 3298 144 3302
rect 148 3298 149 3302
rect 143 3296 149 3298
rect 143 3292 144 3296
rect 148 3292 149 3296
rect 143 3290 149 3292
rect 143 3286 144 3290
rect 148 3286 149 3290
rect 143 3284 149 3286
rect 143 3280 144 3284
rect 148 3280 149 3284
rect 143 3278 149 3280
rect 143 3274 144 3278
rect 148 3274 149 3278
rect 143 3272 149 3274
rect 143 3268 144 3272
rect 148 3268 149 3272
rect 143 3266 149 3268
rect 143 3262 144 3266
rect 148 3262 149 3266
rect 143 3260 149 3262
rect 143 3256 144 3260
rect 148 3256 149 3260
rect 143 3254 149 3256
rect 143 3250 144 3254
rect 148 3250 149 3254
rect 143 3248 149 3250
rect 143 3244 144 3248
rect 148 3244 149 3248
rect 143 3242 149 3244
rect 143 3238 144 3242
rect 148 3238 149 3242
rect 143 3236 149 3238
rect 143 3232 144 3236
rect 148 3232 149 3236
rect 143 3230 149 3232
rect 143 3226 144 3230
rect 148 3226 149 3230
rect 143 3224 149 3226
rect 143 3220 144 3224
rect 148 3220 149 3224
rect 143 3218 149 3220
rect 143 3214 144 3218
rect 148 3214 149 3218
rect 143 3212 149 3214
rect 143 3208 144 3212
rect 148 3208 149 3212
rect 143 3206 149 3208
rect 143 3202 144 3206
rect 148 3202 149 3206
rect 143 3200 149 3202
rect 143 3196 144 3200
rect 148 3196 149 3200
rect 143 3194 149 3196
rect 143 3190 144 3194
rect 148 3190 149 3194
rect 143 3188 149 3190
rect 143 3184 144 3188
rect 148 3184 149 3188
rect 143 3182 149 3184
rect 143 3178 144 3182
rect 148 3178 149 3182
rect 143 3176 149 3178
rect 143 3172 144 3176
rect 148 3172 149 3176
rect 143 3170 149 3172
rect 143 3166 144 3170
rect 148 3166 149 3170
rect 143 3164 149 3166
rect 143 3160 144 3164
rect 148 3160 149 3164
rect 143 3158 149 3160
rect 143 3154 144 3158
rect 148 3154 149 3158
rect 143 3152 149 3154
rect 143 3148 144 3152
rect 148 3148 149 3152
rect 143 3146 149 3148
rect 143 3142 144 3146
rect 148 3142 149 3146
rect 143 3140 149 3142
rect 143 3136 144 3140
rect 148 3136 149 3140
rect 143 3134 149 3136
rect 143 3130 144 3134
rect 148 3130 149 3134
rect 143 3128 149 3130
rect 143 3124 144 3128
rect 148 3124 149 3128
rect 143 3122 149 3124
rect 143 3118 144 3122
rect 148 3118 149 3122
rect 143 3116 149 3118
rect 143 3112 144 3116
rect 148 3112 149 3116
rect 143 3110 149 3112
rect 143 3106 144 3110
rect 148 3106 149 3110
rect 143 3104 149 3106
rect 143 3100 144 3104
rect 148 3100 149 3104
rect 143 3098 149 3100
rect 143 3094 144 3098
rect 148 3094 149 3098
rect 143 3068 149 3094
rect 143 3064 144 3068
rect 148 3064 149 3068
rect 143 3062 149 3064
rect 143 3058 144 3062
rect 148 3058 149 3062
rect 143 3056 149 3058
rect 143 3052 144 3056
rect 148 3052 149 3056
rect 143 3050 149 3052
rect 143 3046 144 3050
rect 148 3046 149 3050
rect 143 3044 149 3046
rect 143 3040 144 3044
rect 148 3040 149 3044
rect 143 3038 149 3040
rect 143 3034 144 3038
rect 148 3034 149 3038
rect 143 3032 149 3034
rect 143 3028 144 3032
rect 148 3028 149 3032
rect 143 3026 149 3028
rect 143 3022 144 3026
rect 148 3022 149 3026
rect 143 3020 149 3022
rect 143 3016 144 3020
rect 148 3016 149 3020
rect 143 3014 149 3016
rect 143 3010 144 3014
rect 148 3010 149 3014
rect 143 3008 149 3010
rect 143 3004 144 3008
rect 148 3004 149 3008
rect 143 3002 149 3004
rect 143 2998 144 3002
rect 148 2998 149 3002
rect 143 2996 149 2998
rect 143 2992 144 2996
rect 148 2992 149 2996
rect 143 2990 149 2992
rect 143 2986 144 2990
rect 148 2986 149 2990
rect 143 2984 149 2986
rect 143 2980 144 2984
rect 148 2980 149 2984
rect 143 2978 149 2980
rect 143 2974 144 2978
rect 148 2974 149 2978
rect 143 2972 149 2974
rect 143 2968 144 2972
rect 148 2968 149 2972
rect 143 2966 149 2968
rect 143 2962 144 2966
rect 148 2962 149 2966
rect 143 2960 149 2962
rect 143 2956 144 2960
rect 148 2956 149 2960
rect 143 2954 149 2956
rect 143 2950 144 2954
rect 148 2950 149 2954
rect 143 2948 149 2950
rect 143 2944 144 2948
rect 148 2944 149 2948
rect 143 2942 149 2944
rect 143 2938 144 2942
rect 148 2938 149 2942
rect 143 2936 149 2938
rect 143 2932 144 2936
rect 148 2932 149 2936
rect 143 2930 149 2932
rect 143 2926 144 2930
rect 148 2926 149 2930
rect 143 2924 149 2926
rect 143 2920 144 2924
rect 148 2920 149 2924
rect 143 2918 149 2920
rect 143 2914 144 2918
rect 148 2914 149 2918
rect 143 2912 149 2914
rect 143 2908 144 2912
rect 148 2908 149 2912
rect 143 2906 149 2908
rect 143 2902 144 2906
rect 148 2902 149 2906
rect 143 2900 149 2902
rect 143 2896 144 2900
rect 148 2896 149 2900
rect 143 2894 149 2896
rect 143 2890 144 2894
rect 148 2890 149 2894
rect 143 2888 149 2890
rect 143 2884 144 2888
rect 148 2884 149 2888
rect 143 2882 149 2884
rect 143 2878 144 2882
rect 148 2878 149 2882
rect 143 2876 149 2878
rect 143 2872 144 2876
rect 148 2872 149 2876
rect 143 2870 149 2872
rect 143 2866 144 2870
rect 148 2866 149 2870
rect 143 2864 149 2866
rect 143 2860 144 2864
rect 148 2860 149 2864
rect 143 2858 149 2860
rect 143 2854 144 2858
rect 148 2854 149 2858
rect 143 2852 149 2854
rect 143 2848 144 2852
rect 148 2848 149 2852
rect 143 2847 149 2848
rect 143 2846 511 2847
rect 143 2842 144 2846
rect 148 2842 150 2846
rect 154 2842 156 2846
rect 160 2842 162 2846
rect 166 2842 168 2846
rect 172 2842 174 2846
rect 178 2842 180 2846
rect 184 2842 186 2846
rect 190 2842 192 2846
rect 196 2842 198 2846
rect 202 2842 204 2846
rect 208 2842 210 2846
rect 214 2842 216 2846
rect 220 2842 222 2846
rect 226 2842 228 2846
rect 232 2842 234 2846
rect 238 2842 240 2846
rect 244 2842 246 2846
rect 250 2842 252 2846
rect 256 2842 258 2846
rect 262 2842 264 2846
rect 268 2842 270 2846
rect 274 2842 276 2846
rect 280 2842 282 2846
rect 286 2842 288 2846
rect 292 2842 294 2846
rect 298 2842 300 2846
rect 304 2842 306 2846
rect 310 2842 312 2846
rect 316 2842 318 2846
rect 322 2842 324 2846
rect 328 2842 330 2846
rect 334 2842 336 2846
rect 340 2842 342 2846
rect 346 2842 348 2846
rect 352 2842 354 2846
rect 358 2842 360 2846
rect 364 2842 366 2846
rect 370 2842 372 2846
rect 376 2842 378 2846
rect 382 2842 384 2846
rect 388 2842 390 2846
rect 394 2842 396 2846
rect 400 2842 402 2846
rect 406 2842 408 2846
rect 412 2842 414 2846
rect 418 2842 420 2846
rect 424 2842 426 2846
rect 430 2842 432 2846
rect 436 2842 438 2846
rect 442 2842 444 2846
rect 448 2842 450 2846
rect 454 2842 456 2846
rect 460 2842 462 2846
rect 466 2842 468 2846
rect 472 2842 474 2846
rect 478 2842 480 2846
rect 484 2842 486 2846
rect 490 2842 492 2846
rect 496 2842 498 2846
rect 502 2842 504 2846
rect 508 2842 511 2846
rect 143 2841 511 2842
rect 143 2840 149 2841
rect 143 2836 144 2840
rect 148 2836 149 2840
rect 143 2834 149 2836
rect 143 2830 144 2834
rect 148 2830 149 2834
rect 143 2828 149 2830
rect 143 2824 144 2828
rect 148 2824 149 2828
rect 143 2822 149 2824
rect 143 2818 144 2822
rect 148 2818 149 2822
rect 143 2816 149 2818
rect 143 2812 144 2816
rect 148 2812 149 2816
rect 143 2810 149 2812
rect 143 2806 144 2810
rect 148 2806 149 2810
rect 143 2804 149 2806
rect 143 2800 144 2804
rect 148 2800 149 2804
rect 143 2798 149 2800
rect 143 2794 144 2798
rect 148 2794 149 2798
rect 143 2792 149 2794
rect 143 2788 144 2792
rect 148 2788 149 2792
rect 143 2786 149 2788
rect 143 2782 144 2786
rect 148 2782 149 2786
rect 143 2780 149 2782
rect 143 2776 144 2780
rect 148 2776 149 2780
rect 143 2774 149 2776
rect 143 2770 144 2774
rect 148 2770 149 2774
rect 143 2768 149 2770
rect 143 2764 144 2768
rect 148 2764 149 2768
rect 143 2762 149 2764
rect 143 2758 144 2762
rect 148 2758 149 2762
rect 143 2756 149 2758
rect 143 2752 144 2756
rect 148 2752 149 2756
rect 143 2750 149 2752
rect 143 2746 144 2750
rect 148 2746 149 2750
rect 143 2744 149 2746
rect 143 2740 144 2744
rect 148 2740 149 2744
rect 143 2738 149 2740
rect 143 2734 144 2738
rect 148 2734 149 2738
rect 143 2732 149 2734
rect 143 2728 144 2732
rect 148 2728 149 2732
rect 143 2726 149 2728
rect 143 2722 144 2726
rect 148 2722 149 2726
rect 143 2720 149 2722
rect 143 2716 144 2720
rect 148 2716 149 2720
rect 143 2714 149 2716
rect 143 2710 144 2714
rect 148 2710 149 2714
rect 143 2708 149 2710
rect 143 2704 144 2708
rect 148 2704 149 2708
rect 143 2702 149 2704
rect 143 2698 144 2702
rect 148 2698 149 2702
rect 143 2696 149 2698
rect 143 2692 144 2696
rect 148 2692 149 2696
rect 143 2690 149 2692
rect 143 2686 144 2690
rect 148 2686 149 2690
rect 143 2684 149 2686
rect 143 2680 144 2684
rect 148 2680 149 2684
rect 143 2678 149 2680
rect 143 2674 144 2678
rect 148 2674 149 2678
rect 143 2672 149 2674
rect 143 2668 144 2672
rect 148 2668 149 2672
rect 143 2666 149 2668
rect 143 2662 144 2666
rect 148 2662 149 2666
rect 143 2660 149 2662
rect 143 2656 144 2660
rect 148 2656 149 2660
rect 143 2654 149 2656
rect 143 2650 144 2654
rect 148 2650 149 2654
rect 143 2648 149 2650
rect 143 2644 144 2648
rect 148 2644 149 2648
rect 143 2642 149 2644
rect 143 2638 144 2642
rect 148 2638 149 2642
rect 143 2636 149 2638
rect 143 2632 144 2636
rect 148 2632 149 2636
rect 143 2630 149 2632
rect 143 2626 144 2630
rect 148 2626 149 2630
rect 143 2624 149 2626
rect 143 2620 144 2624
rect 148 2620 149 2624
rect 143 2594 149 2620
rect 143 2590 144 2594
rect 148 2590 149 2594
rect 143 2588 149 2590
rect 143 2584 144 2588
rect 148 2584 149 2588
rect 143 2582 149 2584
rect 143 2578 144 2582
rect 148 2578 149 2582
rect 143 2576 149 2578
rect 143 2572 144 2576
rect 148 2572 149 2576
rect 143 2570 149 2572
rect 143 2566 144 2570
rect 148 2566 149 2570
rect 143 2564 149 2566
rect 143 2560 144 2564
rect 148 2560 149 2564
rect 143 2558 149 2560
rect 143 2554 144 2558
rect 148 2554 149 2558
rect 143 2552 149 2554
rect 143 2548 144 2552
rect 148 2548 149 2552
rect 143 2546 149 2548
rect 143 2542 144 2546
rect 148 2542 149 2546
rect 143 2540 149 2542
rect 143 2536 144 2540
rect 148 2536 149 2540
rect 143 2534 149 2536
rect 143 2530 144 2534
rect 148 2530 149 2534
rect 143 2528 149 2530
rect 143 2524 144 2528
rect 148 2524 149 2528
rect 143 2522 149 2524
rect 143 2518 144 2522
rect 148 2518 149 2522
rect 143 2516 149 2518
rect 143 2512 144 2516
rect 148 2512 149 2516
rect 143 2510 149 2512
rect 143 2506 144 2510
rect 148 2506 149 2510
rect 143 2504 149 2506
rect 143 2500 144 2504
rect 148 2500 149 2504
rect 143 2498 149 2500
rect 143 2494 144 2498
rect 148 2494 149 2498
rect 143 2492 149 2494
rect 143 2488 144 2492
rect 148 2488 149 2492
rect 143 2486 149 2488
rect 143 2482 144 2486
rect 148 2482 149 2486
rect 143 2480 149 2482
rect 143 2476 144 2480
rect 148 2476 149 2480
rect 143 2474 149 2476
rect 143 2470 144 2474
rect 148 2470 149 2474
rect 143 2468 149 2470
rect 143 2464 144 2468
rect 148 2464 149 2468
rect 143 2462 149 2464
rect 143 2458 144 2462
rect 148 2458 149 2462
rect 143 2456 149 2458
rect 143 2452 144 2456
rect 148 2452 149 2456
rect 143 2450 149 2452
rect 143 2446 144 2450
rect 148 2446 149 2450
rect 143 2444 149 2446
rect 143 2440 144 2444
rect 148 2440 149 2444
rect 143 2438 149 2440
rect 143 2434 144 2438
rect 148 2434 149 2438
rect 143 2432 149 2434
rect 143 2428 144 2432
rect 148 2428 149 2432
rect 143 2426 149 2428
rect 143 2422 144 2426
rect 148 2422 149 2426
rect 143 2420 149 2422
rect 143 2416 144 2420
rect 148 2416 149 2420
rect 143 2414 149 2416
rect 143 2410 144 2414
rect 148 2410 149 2414
rect 143 2408 149 2410
rect 143 2404 144 2408
rect 148 2404 149 2408
rect 143 2402 149 2404
rect 143 2398 144 2402
rect 148 2398 149 2402
rect 143 2396 149 2398
rect 143 2392 144 2396
rect 148 2392 149 2396
rect 143 2390 149 2392
rect 143 2386 144 2390
rect 148 2386 149 2390
rect 143 2384 149 2386
rect 143 2380 144 2384
rect 148 2380 149 2384
rect 143 2378 149 2380
rect 143 2374 144 2378
rect 148 2374 149 2378
rect 143 2373 149 2374
rect 143 2372 511 2373
rect 143 2368 144 2372
rect 148 2368 150 2372
rect 154 2368 156 2372
rect 160 2368 162 2372
rect 166 2368 168 2372
rect 172 2368 174 2372
rect 178 2368 180 2372
rect 184 2368 186 2372
rect 190 2368 192 2372
rect 196 2368 198 2372
rect 202 2368 204 2372
rect 208 2368 210 2372
rect 214 2368 216 2372
rect 220 2368 222 2372
rect 226 2368 228 2372
rect 232 2368 234 2372
rect 238 2368 240 2372
rect 244 2368 246 2372
rect 250 2368 252 2372
rect 256 2368 258 2372
rect 262 2368 264 2372
rect 268 2368 270 2372
rect 274 2368 276 2372
rect 280 2368 282 2372
rect 286 2368 288 2372
rect 292 2368 294 2372
rect 298 2368 300 2372
rect 304 2368 306 2372
rect 310 2368 312 2372
rect 316 2368 318 2372
rect 322 2368 324 2372
rect 328 2368 330 2372
rect 334 2368 336 2372
rect 340 2368 342 2372
rect 346 2368 348 2372
rect 352 2368 354 2372
rect 358 2368 360 2372
rect 364 2368 366 2372
rect 370 2368 372 2372
rect 376 2368 378 2372
rect 382 2368 384 2372
rect 388 2368 390 2372
rect 394 2368 396 2372
rect 400 2368 402 2372
rect 406 2368 408 2372
rect 412 2368 414 2372
rect 418 2368 420 2372
rect 424 2368 426 2372
rect 430 2368 432 2372
rect 436 2368 438 2372
rect 442 2368 444 2372
rect 448 2368 450 2372
rect 454 2368 456 2372
rect 460 2368 462 2372
rect 466 2368 468 2372
rect 472 2368 474 2372
rect 478 2368 480 2372
rect 484 2368 486 2372
rect 490 2368 492 2372
rect 496 2368 498 2372
rect 502 2368 504 2372
rect 508 2368 511 2372
rect 143 2367 511 2368
rect 143 2366 149 2367
rect 143 2362 144 2366
rect 148 2362 149 2366
rect 143 2360 149 2362
rect 143 2356 144 2360
rect 148 2356 149 2360
rect 143 2354 149 2356
rect 143 2350 144 2354
rect 148 2350 149 2354
rect 143 2348 149 2350
rect 143 2344 144 2348
rect 148 2344 149 2348
rect 143 2342 149 2344
rect 143 2338 144 2342
rect 148 2338 149 2342
rect 143 2336 149 2338
rect 143 2332 144 2336
rect 148 2332 149 2336
rect 143 2330 149 2332
rect 143 2326 144 2330
rect 148 2326 149 2330
rect 143 2324 149 2326
rect 143 2320 144 2324
rect 148 2320 149 2324
rect 143 2318 149 2320
rect 143 2314 144 2318
rect 148 2314 149 2318
rect 143 2312 149 2314
rect 143 2308 144 2312
rect 148 2308 149 2312
rect 143 2306 149 2308
rect 143 2302 144 2306
rect 148 2302 149 2306
rect 143 2300 149 2302
rect 143 2296 144 2300
rect 148 2296 149 2300
rect 143 2294 149 2296
rect 143 2290 144 2294
rect 148 2290 149 2294
rect 143 2288 149 2290
rect 143 2284 144 2288
rect 148 2284 149 2288
rect 143 2282 149 2284
rect 143 2278 144 2282
rect 148 2278 149 2282
rect 143 2276 149 2278
rect 143 2272 144 2276
rect 148 2272 149 2276
rect 143 2270 149 2272
rect 143 2266 144 2270
rect 148 2266 149 2270
rect 143 2264 149 2266
rect 143 2260 144 2264
rect 148 2260 149 2264
rect 143 2258 149 2260
rect 143 2254 144 2258
rect 148 2254 149 2258
rect 143 2252 149 2254
rect 143 2248 144 2252
rect 148 2248 149 2252
rect 143 2246 149 2248
rect 143 2242 144 2246
rect 148 2242 149 2246
rect 143 2240 149 2242
rect 143 2236 144 2240
rect 148 2236 149 2240
rect 143 2234 149 2236
rect 143 2230 144 2234
rect 148 2230 149 2234
rect 143 2228 149 2230
rect 143 2224 144 2228
rect 148 2224 149 2228
rect 143 2222 149 2224
rect 143 2218 144 2222
rect 148 2218 149 2222
rect 143 2216 149 2218
rect 143 2212 144 2216
rect 148 2212 149 2216
rect 143 2210 149 2212
rect 143 2206 144 2210
rect 148 2206 149 2210
rect 143 2204 149 2206
rect 143 2200 144 2204
rect 148 2200 149 2204
rect 143 2198 149 2200
rect 143 2194 144 2198
rect 148 2194 149 2198
rect 143 2192 149 2194
rect 143 2188 144 2192
rect 148 2188 149 2192
rect 143 2186 149 2188
rect 143 2182 144 2186
rect 148 2182 149 2186
rect 143 2180 149 2182
rect 143 2176 144 2180
rect 148 2176 149 2180
rect 143 2174 149 2176
rect 143 2170 144 2174
rect 148 2170 149 2174
rect 143 2168 149 2170
rect 143 2164 144 2168
rect 148 2164 149 2168
rect 143 2162 149 2164
rect 143 2158 144 2162
rect 148 2158 149 2162
rect 143 2156 149 2158
rect 143 2152 144 2156
rect 148 2152 149 2156
rect 143 2150 149 2152
rect 143 2146 144 2150
rect 148 2146 149 2150
rect 143 2120 149 2146
rect 143 2116 144 2120
rect 148 2116 149 2120
rect 143 2114 149 2116
rect 143 2110 144 2114
rect 148 2110 149 2114
rect 143 2108 149 2110
rect 143 2104 144 2108
rect 148 2104 149 2108
rect 143 2102 149 2104
rect 143 2098 144 2102
rect 148 2098 149 2102
rect 143 2096 149 2098
rect 143 2092 144 2096
rect 148 2092 149 2096
rect 143 2090 149 2092
rect 143 2086 144 2090
rect 148 2086 149 2090
rect 143 2084 149 2086
rect 143 2080 144 2084
rect 148 2080 149 2084
rect 143 2078 149 2080
rect 143 2074 144 2078
rect 148 2074 149 2078
rect 143 2072 149 2074
rect 143 2068 144 2072
rect 148 2068 149 2072
rect 143 2066 149 2068
rect 143 2062 144 2066
rect 148 2062 149 2066
rect 143 2060 149 2062
rect 143 2056 144 2060
rect 148 2056 149 2060
rect 143 2054 149 2056
rect 143 2050 144 2054
rect 148 2050 149 2054
rect 143 2048 149 2050
rect 143 2044 144 2048
rect 148 2044 149 2048
rect 143 2042 149 2044
rect 143 2038 144 2042
rect 148 2038 149 2042
rect 143 2036 149 2038
rect 143 2032 144 2036
rect 148 2032 149 2036
rect 143 2030 149 2032
rect 143 2026 144 2030
rect 148 2026 149 2030
rect 143 2024 149 2026
rect 143 2020 144 2024
rect 148 2020 149 2024
rect 143 2018 149 2020
rect 143 2014 144 2018
rect 148 2014 149 2018
rect 143 2012 149 2014
rect 143 2008 144 2012
rect 148 2008 149 2012
rect 143 2006 149 2008
rect 143 2002 144 2006
rect 148 2002 149 2006
rect 143 2000 149 2002
rect 143 1996 144 2000
rect 148 1996 149 2000
rect 143 1994 149 1996
rect 143 1990 144 1994
rect 148 1990 149 1994
rect 143 1988 149 1990
rect 143 1984 144 1988
rect 148 1984 149 1988
rect 143 1982 149 1984
rect 143 1978 144 1982
rect 148 1978 149 1982
rect 143 1976 149 1978
rect 143 1972 144 1976
rect 148 1972 149 1976
rect 143 1970 149 1972
rect 143 1966 144 1970
rect 148 1966 149 1970
rect 143 1964 149 1966
rect 143 1960 144 1964
rect 148 1960 149 1964
rect 143 1958 149 1960
rect 143 1954 144 1958
rect 148 1954 149 1958
rect 143 1952 149 1954
rect 143 1948 144 1952
rect 148 1948 149 1952
rect 143 1946 149 1948
rect 143 1942 144 1946
rect 148 1942 149 1946
rect 143 1940 149 1942
rect 143 1936 144 1940
rect 148 1936 149 1940
rect 143 1934 149 1936
rect 143 1930 144 1934
rect 148 1930 149 1934
rect 143 1928 149 1930
rect 143 1924 144 1928
rect 148 1924 149 1928
rect 143 1922 149 1924
rect 143 1918 144 1922
rect 148 1918 149 1922
rect 143 1916 149 1918
rect 143 1912 144 1916
rect 148 1912 149 1916
rect 143 1910 149 1912
rect 143 1906 144 1910
rect 148 1906 149 1910
rect 143 1904 149 1906
rect 143 1900 144 1904
rect 148 1900 149 1904
rect 143 1899 149 1900
rect 143 1898 511 1899
rect 143 1894 144 1898
rect 148 1894 150 1898
rect 154 1894 156 1898
rect 160 1894 162 1898
rect 166 1894 168 1898
rect 172 1894 174 1898
rect 178 1894 180 1898
rect 184 1894 186 1898
rect 190 1894 192 1898
rect 196 1894 198 1898
rect 202 1894 204 1898
rect 208 1894 210 1898
rect 214 1894 216 1898
rect 220 1894 222 1898
rect 226 1894 228 1898
rect 232 1894 234 1898
rect 238 1894 240 1898
rect 244 1894 246 1898
rect 250 1894 252 1898
rect 256 1894 258 1898
rect 262 1894 264 1898
rect 268 1894 270 1898
rect 274 1894 276 1898
rect 280 1894 282 1898
rect 286 1894 288 1898
rect 292 1894 294 1898
rect 298 1894 300 1898
rect 304 1894 306 1898
rect 310 1894 312 1898
rect 316 1894 318 1898
rect 322 1894 324 1898
rect 328 1894 330 1898
rect 334 1894 336 1898
rect 340 1894 342 1898
rect 346 1894 348 1898
rect 352 1894 354 1898
rect 358 1894 360 1898
rect 364 1894 366 1898
rect 370 1894 372 1898
rect 376 1894 378 1898
rect 382 1894 384 1898
rect 388 1894 390 1898
rect 394 1894 396 1898
rect 400 1894 402 1898
rect 406 1894 408 1898
rect 412 1894 414 1898
rect 418 1894 420 1898
rect 424 1894 426 1898
rect 430 1894 432 1898
rect 436 1894 438 1898
rect 442 1894 444 1898
rect 448 1894 450 1898
rect 454 1894 456 1898
rect 460 1894 462 1898
rect 466 1894 468 1898
rect 472 1894 474 1898
rect 478 1894 480 1898
rect 484 1894 486 1898
rect 490 1894 492 1898
rect 496 1894 498 1898
rect 502 1894 504 1898
rect 508 1894 511 1898
rect 143 1893 511 1894
rect 143 1892 149 1893
rect 143 1888 144 1892
rect 148 1888 149 1892
rect 143 1886 149 1888
rect 143 1882 144 1886
rect 148 1882 149 1886
rect 143 1880 149 1882
rect 143 1876 144 1880
rect 148 1876 149 1880
rect 143 1874 149 1876
rect 143 1870 144 1874
rect 148 1870 149 1874
rect 143 1868 149 1870
rect 143 1864 144 1868
rect 148 1864 149 1868
rect 143 1862 149 1864
rect 143 1858 144 1862
rect 148 1858 149 1862
rect 143 1856 149 1858
rect 143 1852 144 1856
rect 148 1852 149 1856
rect 143 1850 149 1852
rect 143 1846 144 1850
rect 148 1846 149 1850
rect 143 1844 149 1846
rect 143 1840 144 1844
rect 148 1840 149 1844
rect 143 1838 149 1840
rect 143 1834 144 1838
rect 148 1834 149 1838
rect 143 1832 149 1834
rect 143 1828 144 1832
rect 148 1828 149 1832
rect 143 1826 149 1828
rect 143 1822 144 1826
rect 148 1822 149 1826
rect 143 1820 149 1822
rect 143 1816 144 1820
rect 148 1816 149 1820
rect 143 1814 149 1816
rect 143 1810 144 1814
rect 148 1810 149 1814
rect 143 1808 149 1810
rect 143 1804 144 1808
rect 148 1804 149 1808
rect 143 1802 149 1804
rect 143 1798 144 1802
rect 148 1798 149 1802
rect 143 1796 149 1798
rect 143 1792 144 1796
rect 148 1792 149 1796
rect 143 1790 149 1792
rect 143 1786 144 1790
rect 148 1786 149 1790
rect 143 1784 149 1786
rect 143 1780 144 1784
rect 148 1780 149 1784
rect 143 1778 149 1780
rect 143 1774 144 1778
rect 148 1774 149 1778
rect 143 1772 149 1774
rect 143 1768 144 1772
rect 148 1768 149 1772
rect 143 1766 149 1768
rect 143 1762 144 1766
rect 148 1762 149 1766
rect 143 1760 149 1762
rect 143 1756 144 1760
rect 148 1756 149 1760
rect 143 1754 149 1756
rect 143 1750 144 1754
rect 148 1750 149 1754
rect 143 1748 149 1750
rect 143 1744 144 1748
rect 148 1744 149 1748
rect 143 1742 149 1744
rect 143 1738 144 1742
rect 148 1738 149 1742
rect 143 1736 149 1738
rect 143 1732 144 1736
rect 148 1732 149 1736
rect 143 1730 149 1732
rect 143 1726 144 1730
rect 148 1726 149 1730
rect 143 1724 149 1726
rect 143 1720 144 1724
rect 148 1720 149 1724
rect 143 1718 149 1720
rect 143 1714 144 1718
rect 148 1714 149 1718
rect 143 1712 149 1714
rect 143 1708 144 1712
rect 148 1708 149 1712
rect 143 1706 149 1708
rect 143 1702 144 1706
rect 148 1702 149 1706
rect 143 1700 149 1702
rect 143 1696 144 1700
rect 148 1696 149 1700
rect 143 1694 149 1696
rect 143 1690 144 1694
rect 148 1690 149 1694
rect 143 1688 149 1690
rect 143 1684 144 1688
rect 148 1684 149 1688
rect 143 1682 149 1684
rect 143 1678 144 1682
rect 148 1678 149 1682
rect 143 1676 149 1678
rect 143 1672 144 1676
rect 148 1672 149 1676
rect 143 1646 149 1672
rect 143 1642 144 1646
rect 148 1642 149 1646
rect 143 1640 149 1642
rect 143 1636 144 1640
rect 148 1636 149 1640
rect 143 1634 149 1636
rect 143 1630 144 1634
rect 148 1630 149 1634
rect 143 1628 149 1630
rect 143 1624 144 1628
rect 148 1624 149 1628
rect 143 1622 149 1624
rect 143 1618 144 1622
rect 148 1618 149 1622
rect 143 1616 149 1618
rect 143 1612 144 1616
rect 148 1612 149 1616
rect 143 1610 149 1612
rect 143 1606 144 1610
rect 148 1606 149 1610
rect 143 1604 149 1606
rect 143 1600 144 1604
rect 148 1600 149 1604
rect 143 1598 149 1600
rect 143 1594 144 1598
rect 148 1594 149 1598
rect 143 1592 149 1594
rect 143 1588 144 1592
rect 148 1588 149 1592
rect 143 1586 149 1588
rect 143 1582 144 1586
rect 148 1582 149 1586
rect 143 1580 149 1582
rect 143 1576 144 1580
rect 148 1576 149 1580
rect 143 1574 149 1576
rect 143 1570 144 1574
rect 148 1570 149 1574
rect 143 1568 149 1570
rect 143 1564 144 1568
rect 148 1564 149 1568
rect 143 1562 149 1564
rect 143 1558 144 1562
rect 148 1558 149 1562
rect 143 1556 149 1558
rect 143 1552 144 1556
rect 148 1552 149 1556
rect 143 1550 149 1552
rect 143 1546 144 1550
rect 148 1546 149 1550
rect 143 1544 149 1546
rect 143 1540 144 1544
rect 148 1540 149 1544
rect 143 1538 149 1540
rect 143 1534 144 1538
rect 148 1534 149 1538
rect 143 1532 149 1534
rect 143 1528 144 1532
rect 148 1528 149 1532
rect 143 1526 149 1528
rect 143 1522 144 1526
rect 148 1522 149 1526
rect 143 1520 149 1522
rect 143 1516 144 1520
rect 148 1516 149 1520
rect 143 1514 149 1516
rect 143 1510 144 1514
rect 148 1510 149 1514
rect 143 1508 149 1510
rect 143 1504 144 1508
rect 148 1504 149 1508
rect 143 1502 149 1504
rect 143 1498 144 1502
rect 148 1498 149 1502
rect 143 1496 149 1498
rect 143 1492 144 1496
rect 148 1492 149 1496
rect 143 1490 149 1492
rect 143 1486 144 1490
rect 148 1486 149 1490
rect 143 1484 149 1486
rect 143 1480 144 1484
rect 148 1480 149 1484
rect 143 1478 149 1480
rect 143 1474 144 1478
rect 148 1474 149 1478
rect 143 1472 149 1474
rect 143 1468 144 1472
rect 148 1468 149 1472
rect 143 1466 149 1468
rect 143 1462 144 1466
rect 148 1462 149 1466
rect 143 1460 149 1462
rect 143 1456 144 1460
rect 148 1456 149 1460
rect 143 1454 149 1456
rect 143 1450 144 1454
rect 148 1450 149 1454
rect 143 1448 149 1450
rect 143 1444 144 1448
rect 148 1444 149 1448
rect 143 1442 149 1444
rect 143 1438 144 1442
rect 148 1438 149 1442
rect 143 1436 149 1438
rect 143 1432 144 1436
rect 148 1432 149 1436
rect 143 1430 149 1432
rect 143 1426 144 1430
rect 148 1426 149 1430
rect 143 1425 149 1426
rect 143 1424 511 1425
rect 143 1420 144 1424
rect 148 1420 150 1424
rect 154 1420 156 1424
rect 160 1420 162 1424
rect 166 1420 168 1424
rect 172 1420 174 1424
rect 178 1420 180 1424
rect 184 1420 186 1424
rect 190 1420 192 1424
rect 196 1420 198 1424
rect 202 1420 204 1424
rect 208 1420 210 1424
rect 214 1420 216 1424
rect 220 1420 222 1424
rect 226 1420 228 1424
rect 232 1420 234 1424
rect 238 1420 240 1424
rect 244 1420 246 1424
rect 250 1420 252 1424
rect 256 1420 258 1424
rect 262 1420 264 1424
rect 268 1420 270 1424
rect 274 1420 276 1424
rect 280 1420 282 1424
rect 286 1420 288 1424
rect 292 1420 294 1424
rect 298 1420 300 1424
rect 304 1420 306 1424
rect 310 1420 312 1424
rect 316 1420 318 1424
rect 322 1420 324 1424
rect 328 1420 330 1424
rect 334 1420 336 1424
rect 340 1420 342 1424
rect 346 1420 348 1424
rect 352 1420 354 1424
rect 358 1420 360 1424
rect 364 1420 366 1424
rect 370 1420 372 1424
rect 376 1420 378 1424
rect 382 1420 384 1424
rect 388 1420 390 1424
rect 394 1420 396 1424
rect 400 1420 402 1424
rect 406 1420 408 1424
rect 412 1420 414 1424
rect 418 1420 420 1424
rect 424 1420 426 1424
rect 430 1420 432 1424
rect 436 1420 438 1424
rect 442 1420 444 1424
rect 448 1420 450 1424
rect 454 1420 456 1424
rect 460 1420 462 1424
rect 466 1420 468 1424
rect 472 1420 474 1424
rect 478 1420 480 1424
rect 484 1420 486 1424
rect 490 1420 492 1424
rect 496 1420 498 1424
rect 502 1420 504 1424
rect 508 1420 511 1424
rect 143 1419 511 1420
rect 143 1418 149 1419
rect 143 1414 144 1418
rect 148 1414 149 1418
rect 143 1412 149 1414
rect 143 1408 144 1412
rect 148 1408 149 1412
rect 143 1406 149 1408
rect 143 1402 144 1406
rect 148 1402 149 1406
rect 143 1400 149 1402
rect 143 1396 144 1400
rect 148 1396 149 1400
rect 143 1394 149 1396
rect 143 1390 144 1394
rect 148 1390 149 1394
rect 143 1388 149 1390
rect 143 1384 144 1388
rect 148 1384 149 1388
rect 143 1382 149 1384
rect 143 1378 144 1382
rect 148 1378 149 1382
rect 143 1376 149 1378
rect 143 1372 144 1376
rect 148 1372 149 1376
rect 143 1370 149 1372
rect 143 1366 144 1370
rect 148 1366 149 1370
rect 143 1364 149 1366
rect 143 1360 144 1364
rect 148 1360 149 1364
rect 143 1358 149 1360
rect 143 1354 144 1358
rect 148 1354 149 1358
rect 143 1352 149 1354
rect 143 1348 144 1352
rect 148 1348 149 1352
rect 143 1346 149 1348
rect 143 1342 144 1346
rect 148 1342 149 1346
rect 143 1340 149 1342
rect 143 1336 144 1340
rect 148 1336 149 1340
rect 143 1334 149 1336
rect 143 1330 144 1334
rect 148 1330 149 1334
rect 143 1328 149 1330
rect 143 1324 144 1328
rect 148 1324 149 1328
rect 143 1322 149 1324
rect 143 1318 144 1322
rect 148 1318 149 1322
rect 143 1316 149 1318
rect 143 1312 144 1316
rect 148 1312 149 1316
rect 143 1310 149 1312
rect 143 1306 144 1310
rect 148 1306 149 1310
rect 143 1304 149 1306
rect 143 1300 144 1304
rect 148 1300 149 1304
rect 143 1298 149 1300
rect 143 1294 144 1298
rect 148 1294 149 1298
rect 143 1292 149 1294
rect 143 1288 144 1292
rect 148 1288 149 1292
rect 143 1286 149 1288
rect 143 1282 144 1286
rect 148 1282 149 1286
rect 143 1280 149 1282
rect 143 1276 144 1280
rect 148 1276 149 1280
rect 143 1274 149 1276
rect 143 1270 144 1274
rect 148 1270 149 1274
rect 143 1268 149 1270
rect 143 1264 144 1268
rect 148 1264 149 1268
rect 143 1262 149 1264
rect 143 1258 144 1262
rect 148 1258 149 1262
rect 143 1256 149 1258
rect 143 1252 144 1256
rect 148 1252 149 1256
rect 143 1250 149 1252
rect 143 1246 144 1250
rect 148 1246 149 1250
rect 143 1244 149 1246
rect 143 1240 144 1244
rect 148 1240 149 1244
rect 143 1238 149 1240
rect 143 1234 144 1238
rect 148 1234 149 1238
rect 143 1232 149 1234
rect 143 1228 144 1232
rect 148 1228 149 1232
rect 143 1226 149 1228
rect 143 1222 144 1226
rect 148 1222 149 1226
rect 143 1220 149 1222
rect 143 1216 144 1220
rect 148 1216 149 1220
rect 143 1214 149 1216
rect 143 1210 144 1214
rect 148 1210 149 1214
rect 143 1208 149 1210
rect 143 1204 144 1208
rect 148 1204 149 1208
rect 143 1202 149 1204
rect 143 1198 144 1202
rect 148 1198 149 1202
rect 143 1172 149 1198
rect 143 1168 144 1172
rect 148 1168 149 1172
rect 143 1166 149 1168
rect 143 1162 144 1166
rect 148 1162 149 1166
rect 143 1160 149 1162
rect 143 1156 144 1160
rect 148 1156 149 1160
rect 143 1154 149 1156
rect 143 1150 144 1154
rect 148 1150 149 1154
rect 143 1148 149 1150
rect 143 1144 144 1148
rect 148 1144 149 1148
rect 143 1142 149 1144
rect 143 1138 144 1142
rect 148 1138 149 1142
rect 143 1136 149 1138
rect 143 1132 144 1136
rect 148 1132 149 1136
rect 143 1130 149 1132
rect 143 1126 144 1130
rect 148 1126 149 1130
rect 143 1124 149 1126
rect 143 1120 144 1124
rect 148 1120 149 1124
rect 143 1118 149 1120
rect 143 1114 144 1118
rect 148 1114 149 1118
rect 143 1112 149 1114
rect 143 1108 144 1112
rect 148 1108 149 1112
rect 143 1106 149 1108
rect 143 1102 144 1106
rect 148 1102 149 1106
rect 143 1100 149 1102
rect 143 1096 144 1100
rect 148 1096 149 1100
rect 143 1094 149 1096
rect 143 1090 144 1094
rect 148 1090 149 1094
rect 143 1088 149 1090
rect 143 1084 144 1088
rect 148 1084 149 1088
rect 143 1082 149 1084
rect 143 1078 144 1082
rect 148 1078 149 1082
rect 143 1076 149 1078
rect 143 1072 144 1076
rect 148 1072 149 1076
rect 143 1070 149 1072
rect 143 1066 144 1070
rect 148 1066 149 1070
rect 143 1064 149 1066
rect 143 1060 144 1064
rect 148 1060 149 1064
rect 143 1058 149 1060
rect 143 1054 144 1058
rect 148 1054 149 1058
rect 143 1052 149 1054
rect 143 1048 144 1052
rect 148 1048 149 1052
rect 143 1046 149 1048
rect 143 1042 144 1046
rect 148 1042 149 1046
rect 143 1040 149 1042
rect 143 1036 144 1040
rect 148 1036 149 1040
rect 143 1034 149 1036
rect 143 1030 144 1034
rect 148 1030 149 1034
rect 143 1028 149 1030
rect 143 1024 144 1028
rect 148 1024 149 1028
rect 143 1022 149 1024
rect 143 1018 144 1022
rect 148 1018 149 1022
rect 143 1016 149 1018
rect 143 1012 144 1016
rect 148 1012 149 1016
rect 143 1010 149 1012
rect 143 1006 144 1010
rect 148 1006 149 1010
rect 143 1004 149 1006
rect 143 1000 144 1004
rect 148 1000 149 1004
rect 143 998 149 1000
rect 143 994 144 998
rect 148 994 149 998
rect 143 992 149 994
rect 143 988 144 992
rect 148 988 149 992
rect 143 986 149 988
rect 143 982 144 986
rect 148 982 149 986
rect 143 980 149 982
rect 143 976 144 980
rect 148 976 149 980
rect 143 974 149 976
rect 143 970 144 974
rect 148 970 149 974
rect 143 968 149 970
rect 143 964 144 968
rect 148 964 149 968
rect 143 962 149 964
rect 143 958 144 962
rect 148 958 149 962
rect 143 956 149 958
rect 143 952 144 956
rect 148 952 149 956
rect 143 951 149 952
rect 143 950 511 951
rect 143 946 144 950
rect 148 946 150 950
rect 154 946 156 950
rect 160 946 162 950
rect 166 946 168 950
rect 172 946 174 950
rect 178 946 180 950
rect 184 946 186 950
rect 190 946 192 950
rect 196 946 198 950
rect 202 946 204 950
rect 208 946 210 950
rect 214 946 216 950
rect 220 946 222 950
rect 226 946 228 950
rect 232 946 234 950
rect 238 946 240 950
rect 244 946 246 950
rect 250 946 252 950
rect 256 946 258 950
rect 262 946 264 950
rect 268 946 270 950
rect 274 946 276 950
rect 280 946 282 950
rect 286 946 288 950
rect 292 946 294 950
rect 298 946 300 950
rect 304 946 306 950
rect 310 946 312 950
rect 316 946 318 950
rect 322 946 324 950
rect 328 946 330 950
rect 334 946 336 950
rect 340 946 342 950
rect 346 946 348 950
rect 352 946 354 950
rect 358 946 360 950
rect 364 946 366 950
rect 370 946 372 950
rect 376 946 378 950
rect 382 946 384 950
rect 388 946 390 950
rect 394 946 396 950
rect 400 946 402 950
rect 406 946 408 950
rect 412 946 414 950
rect 418 946 420 950
rect 424 946 426 950
rect 430 946 432 950
rect 436 946 438 950
rect 442 946 444 950
rect 448 946 450 950
rect 454 946 456 950
rect 460 946 462 950
rect 466 946 468 950
rect 472 946 474 950
rect 478 946 480 950
rect 484 946 486 950
rect 490 946 492 950
rect 496 946 498 950
rect 502 946 504 950
rect 508 946 511 950
rect 143 945 511 946
rect 143 944 149 945
rect 143 940 144 944
rect 148 940 149 944
rect 143 938 149 940
rect 143 934 144 938
rect 148 934 149 938
rect 143 932 149 934
rect 143 928 144 932
rect 148 928 149 932
rect 143 926 149 928
rect 143 922 144 926
rect 148 922 149 926
rect 143 920 149 922
rect 143 916 144 920
rect 148 916 149 920
rect 143 914 149 916
rect 143 910 144 914
rect 148 910 149 914
rect 143 908 149 910
rect 143 904 144 908
rect 148 904 149 908
rect 143 902 149 904
rect 143 898 144 902
rect 148 898 149 902
rect 143 896 149 898
rect 143 892 144 896
rect 148 892 149 896
rect 143 890 149 892
rect 143 886 144 890
rect 148 886 149 890
rect 143 884 149 886
rect 143 880 144 884
rect 148 880 149 884
rect 143 878 149 880
rect 143 874 144 878
rect 148 874 149 878
rect 143 872 149 874
rect 143 868 144 872
rect 148 868 149 872
rect 143 866 149 868
rect 143 862 144 866
rect 148 862 149 866
rect 143 860 149 862
rect 143 856 144 860
rect 148 856 149 860
rect 143 854 149 856
rect 143 850 144 854
rect 148 850 149 854
rect 143 848 149 850
rect 143 844 144 848
rect 148 844 149 848
rect 143 842 149 844
rect 143 838 144 842
rect 148 838 149 842
rect 143 836 149 838
rect 143 832 144 836
rect 148 832 149 836
rect 143 830 149 832
rect 143 826 144 830
rect 148 826 149 830
rect 143 824 149 826
rect 143 820 144 824
rect 148 820 149 824
rect 143 818 149 820
rect 143 814 144 818
rect 148 814 149 818
rect 143 812 149 814
rect 143 808 144 812
rect 148 808 149 812
rect 143 806 149 808
rect 143 802 144 806
rect 148 802 149 806
rect 143 800 149 802
rect 143 796 144 800
rect 148 796 149 800
rect 143 794 149 796
rect 143 790 144 794
rect 148 790 149 794
rect 143 788 149 790
rect 143 784 144 788
rect 148 784 149 788
rect 143 782 149 784
rect 143 778 144 782
rect 148 778 149 782
rect 143 776 149 778
rect 143 772 144 776
rect 148 772 149 776
rect 143 770 149 772
rect 143 766 144 770
rect 148 766 149 770
rect 143 764 149 766
rect 143 760 144 764
rect 148 760 149 764
rect 143 758 149 760
rect 143 754 144 758
rect 148 754 149 758
rect 143 752 149 754
rect 143 748 144 752
rect 148 748 149 752
rect 143 746 149 748
rect 143 742 144 746
rect 148 742 149 746
rect 143 740 149 742
rect 143 736 144 740
rect 148 736 149 740
rect 143 734 149 736
rect 143 730 144 734
rect 148 730 149 734
rect 143 728 149 730
rect 143 724 144 728
rect 148 724 149 728
rect 143 698 149 724
rect 143 694 144 698
rect 148 694 149 698
rect 143 692 149 694
rect 143 688 144 692
rect 148 688 149 692
rect 143 686 149 688
rect 143 682 144 686
rect 148 682 149 686
rect 143 680 149 682
rect 143 676 144 680
rect 148 676 149 680
rect 143 674 149 676
rect 143 670 144 674
rect 148 670 149 674
rect 143 668 149 670
rect 143 664 144 668
rect 148 664 149 668
rect 143 662 149 664
rect 143 658 144 662
rect 148 658 149 662
rect 143 656 149 658
rect 143 652 144 656
rect 148 652 149 656
rect 143 650 149 652
rect 143 646 144 650
rect 148 646 149 650
rect 143 644 149 646
rect 143 640 144 644
rect 148 640 149 644
rect 143 638 149 640
rect 143 634 144 638
rect 148 634 149 638
rect 143 632 149 634
rect 143 628 144 632
rect 148 628 149 632
rect 143 626 149 628
rect 143 622 144 626
rect 148 622 149 626
rect 143 620 149 622
rect 143 616 144 620
rect 148 616 149 620
rect 143 614 149 616
rect 143 610 144 614
rect 148 610 149 614
rect 143 608 149 610
rect 143 604 144 608
rect 148 604 149 608
rect 143 602 149 604
rect 143 598 144 602
rect 148 598 149 602
rect 143 596 149 598
rect 143 592 144 596
rect 148 592 149 596
rect 143 590 149 592
rect 143 586 144 590
rect 148 586 149 590
rect 143 584 149 586
rect 143 580 144 584
rect 148 580 149 584
rect 143 578 149 580
rect 143 574 144 578
rect 148 574 149 578
rect 143 572 149 574
rect 143 568 144 572
rect 148 568 149 572
rect 143 566 149 568
rect 143 562 144 566
rect 148 562 149 566
rect 143 560 149 562
rect 143 556 144 560
rect 148 556 149 560
rect 143 554 149 556
rect 143 550 144 554
rect 148 550 149 554
rect 143 548 149 550
rect 143 544 144 548
rect 148 544 149 548
rect 143 542 149 544
rect 143 538 144 542
rect 148 538 149 542
rect 143 536 149 538
rect 143 532 144 536
rect 148 532 149 536
rect 143 530 149 532
rect 143 526 144 530
rect 148 526 149 530
rect 143 524 149 526
rect 143 520 144 524
rect 148 520 149 524
rect 143 518 149 520
rect 143 514 144 518
rect 148 514 149 518
rect 143 512 149 514
rect 143 508 144 512
rect 148 508 149 512
rect 143 506 149 508
rect 143 502 144 506
rect 148 502 149 506
rect 143 500 149 502
rect 143 496 144 500
rect 148 496 149 500
rect 143 494 149 496
rect 143 490 144 494
rect 148 490 149 494
rect 143 488 149 490
rect 143 484 144 488
rect 148 484 149 488
rect 143 482 149 484
rect 143 478 144 482
rect 148 478 149 482
rect 143 477 149 478
rect 143 476 511 477
rect 143 472 144 476
rect 148 472 150 476
rect 154 472 156 476
rect 160 472 162 476
rect 166 472 168 476
rect 172 472 174 476
rect 178 472 180 476
rect 184 472 186 476
rect 190 472 192 476
rect 196 472 198 476
rect 202 472 204 476
rect 208 472 210 476
rect 214 472 216 476
rect 220 472 222 476
rect 226 472 228 476
rect 232 472 234 476
rect 238 472 240 476
rect 244 472 246 476
rect 250 472 252 476
rect 256 472 258 476
rect 262 472 264 476
rect 268 472 270 476
rect 274 472 276 476
rect 280 472 282 476
rect 286 472 288 476
rect 292 472 294 476
rect 298 472 300 476
rect 304 472 306 476
rect 310 472 312 476
rect 316 472 318 476
rect 322 472 324 476
rect 328 472 330 476
rect 334 472 336 476
rect 340 472 342 476
rect 346 472 348 476
rect 352 472 354 476
rect 358 472 360 476
rect 364 472 366 476
rect 370 472 372 476
rect 376 472 378 476
rect 382 472 384 476
rect 388 472 390 476
rect 394 472 396 476
rect 400 472 402 476
rect 406 472 408 476
rect 412 472 414 476
rect 418 472 420 476
rect 424 472 426 476
rect 430 472 432 476
rect 436 472 438 476
rect 442 472 444 476
rect 448 472 450 476
rect 454 472 456 476
rect 460 472 462 476
rect 466 472 468 476
rect 472 472 474 476
rect 478 472 480 476
rect 484 472 486 476
rect 490 472 492 476
rect 496 472 498 476
rect 502 472 504 476
rect 508 472 511 476
rect 143 471 511 472
rect 143 470 149 471
rect 143 466 144 470
rect 148 466 149 470
rect 143 464 149 466
rect 143 460 144 464
rect 148 460 149 464
rect 143 458 149 460
rect 143 454 144 458
rect 148 454 149 458
rect 143 452 149 454
rect 143 448 144 452
rect 148 448 149 452
rect 143 446 149 448
rect 143 442 144 446
rect 148 442 149 446
rect 143 440 149 442
rect 143 436 144 440
rect 148 436 149 440
rect 143 434 149 436
rect 143 430 144 434
rect 148 430 149 434
rect 143 428 149 430
rect 143 424 144 428
rect 148 424 149 428
rect 143 422 149 424
rect 143 418 144 422
rect 148 418 149 422
rect 143 416 149 418
rect 143 412 144 416
rect 148 412 149 416
rect 143 410 149 412
rect 143 406 144 410
rect 148 406 149 410
rect 143 404 149 406
rect 143 400 144 404
rect 148 400 149 404
rect 143 398 149 400
rect 143 394 144 398
rect 148 394 149 398
rect 143 392 149 394
rect 143 388 144 392
rect 148 388 149 392
rect 143 386 149 388
rect 143 382 144 386
rect 148 382 149 386
rect 143 380 149 382
rect 143 376 144 380
rect 148 376 149 380
rect 143 374 149 376
rect 143 370 144 374
rect 148 370 149 374
rect 143 368 149 370
rect 143 364 144 368
rect 148 364 149 368
rect 143 362 149 364
rect 143 358 144 362
rect 148 358 149 362
rect 143 356 149 358
rect 143 352 144 356
rect 148 352 149 356
rect 143 350 149 352
rect 143 346 144 350
rect 148 346 149 350
rect 143 344 149 346
rect 143 340 144 344
rect 148 340 149 344
rect 143 338 149 340
rect 143 334 144 338
rect 148 334 149 338
rect 143 332 149 334
rect 143 328 144 332
rect 148 328 149 332
rect 143 326 149 328
rect 143 322 144 326
rect 148 322 149 326
rect 143 320 149 322
rect 143 316 144 320
rect 148 316 149 320
rect 143 314 149 316
rect 143 310 144 314
rect 148 310 149 314
rect 143 308 149 310
rect 143 304 144 308
rect 148 304 149 308
rect 143 302 149 304
rect 143 298 144 302
rect 148 298 149 302
rect 143 296 149 298
rect 143 292 144 296
rect 148 292 149 296
rect 143 290 149 292
rect 143 286 144 290
rect 148 286 149 290
rect 143 284 149 286
rect 143 280 144 284
rect 148 280 149 284
rect 143 278 149 280
rect 143 274 144 278
rect 148 274 149 278
rect 143 272 149 274
rect 143 268 144 272
rect 148 268 149 272
rect 143 266 149 268
rect 143 262 144 266
rect 148 262 149 266
rect 143 260 149 262
rect 143 256 144 260
rect 148 256 149 260
rect 143 254 149 256
rect 143 250 144 254
rect 148 250 149 254
rect 143 224 149 250
rect 143 220 144 224
rect 148 220 149 224
rect 143 218 149 220
rect 143 214 144 218
rect 148 214 149 218
rect 143 212 149 214
rect 143 208 144 212
rect 148 208 149 212
rect 143 206 149 208
rect 143 202 144 206
rect 148 202 149 206
rect 143 200 149 202
rect 143 196 144 200
rect 148 196 149 200
rect 143 194 149 196
rect 143 190 144 194
rect 148 190 149 194
rect 143 188 149 190
rect 143 184 144 188
rect 148 184 149 188
rect 143 182 149 184
rect 143 178 144 182
rect 148 178 149 182
rect 143 176 149 178
rect 143 172 144 176
rect 148 172 149 176
rect 143 170 149 172
rect 143 166 144 170
rect 148 166 149 170
rect 143 164 149 166
rect 143 160 144 164
rect 148 160 149 164
rect 143 158 149 160
rect 143 154 144 158
rect 148 154 149 158
rect 143 152 149 154
rect 143 148 144 152
rect 148 148 149 152
rect 143 146 149 148
rect 143 142 144 146
rect 148 142 149 146
rect 143 140 149 142
rect 143 136 144 140
rect 148 136 149 140
rect 143 134 149 136
rect 143 130 144 134
rect 148 130 149 134
rect 143 128 149 130
rect 143 124 144 128
rect 148 124 149 128
rect 143 122 149 124
rect 143 118 144 122
rect 148 118 149 122
rect 143 116 149 118
rect 143 112 144 116
rect 148 112 149 116
rect 143 110 149 112
rect 143 106 144 110
rect 148 106 149 110
rect 143 104 149 106
rect 143 100 144 104
rect 148 100 149 104
rect 143 98 149 100
rect 143 94 144 98
rect 148 94 149 98
rect 143 92 149 94
rect 143 88 144 92
rect 148 88 149 92
rect 143 86 149 88
rect 143 82 144 86
rect 148 82 149 86
rect 143 80 149 82
rect 143 76 144 80
rect 148 76 149 80
rect 143 74 149 76
rect 143 70 144 74
rect 148 70 149 74
rect 143 68 149 70
rect 143 64 144 68
rect 148 64 149 68
rect 143 62 149 64
rect 143 58 144 62
rect 148 58 149 62
rect 143 56 149 58
rect 143 52 144 56
rect 148 52 149 56
rect 143 50 149 52
rect 143 46 144 50
rect 148 46 149 50
rect 143 44 149 46
rect 143 40 144 44
rect 148 40 149 44
rect 143 38 149 40
rect 143 34 144 38
rect 148 34 149 38
rect 143 32 149 34
rect 143 28 144 32
rect 148 28 149 32
rect 143 26 149 28
rect 143 22 144 26
rect 148 22 149 26
rect 143 20 149 22
rect 143 16 144 20
rect 148 16 149 20
rect 143 14 149 16
rect 143 10 144 14
rect 148 10 149 14
rect 143 8 149 10
rect 143 4 144 8
rect 148 4 149 8
rect 143 3 149 4
<< psubstratepcontact >>
rect 144 4258 148 4262
rect 144 4252 148 4256
rect 144 4246 148 4250
rect 144 4240 148 4244
rect 144 4234 148 4238
rect 144 4228 148 4232
rect 144 4222 148 4226
rect 144 4216 148 4220
rect 144 4210 148 4214
rect 144 4204 148 4208
rect 144 4198 148 4202
rect 144 4192 148 4196
rect 144 4186 148 4190
rect 144 4180 148 4184
rect 144 4174 148 4178
rect 144 4168 148 4172
rect 144 4162 148 4166
rect 144 4156 148 4160
rect 144 4150 148 4154
rect 144 4144 148 4148
rect 144 4138 148 4142
rect 144 4132 148 4136
rect 144 4126 148 4130
rect 144 4120 148 4124
rect 144 4114 148 4118
rect 144 4108 148 4112
rect 144 4102 148 4106
rect 144 4096 148 4100
rect 144 4090 148 4094
rect 144 4084 148 4088
rect 144 4078 148 4082
rect 144 4072 148 4076
rect 144 4066 148 4070
rect 144 4060 148 4064
rect 144 4054 148 4058
rect 144 4048 148 4052
rect 144 4042 148 4046
rect 144 4012 148 4016
rect 144 4006 148 4010
rect 144 4000 148 4004
rect 144 3994 148 3998
rect 144 3988 148 3992
rect 144 3982 148 3986
rect 144 3976 148 3980
rect 144 3970 148 3974
rect 144 3964 148 3968
rect 144 3958 148 3962
rect 144 3952 148 3956
rect 144 3946 148 3950
rect 144 3940 148 3944
rect 144 3934 148 3938
rect 144 3928 148 3932
rect 144 3922 148 3926
rect 144 3916 148 3920
rect 144 3910 148 3914
rect 144 3904 148 3908
rect 144 3898 148 3902
rect 144 3892 148 3896
rect 144 3886 148 3890
rect 144 3880 148 3884
rect 144 3874 148 3878
rect 144 3868 148 3872
rect 144 3862 148 3866
rect 144 3856 148 3860
rect 144 3850 148 3854
rect 144 3844 148 3848
rect 144 3838 148 3842
rect 144 3832 148 3836
rect 144 3826 148 3830
rect 144 3820 148 3824
rect 144 3814 148 3818
rect 144 3808 148 3812
rect 144 3802 148 3806
rect 144 3796 148 3800
rect 144 3790 148 3794
rect 150 3790 154 3794
rect 156 3790 160 3794
rect 162 3790 166 3794
rect 168 3790 172 3794
rect 174 3790 178 3794
rect 180 3790 184 3794
rect 186 3790 190 3794
rect 192 3790 196 3794
rect 198 3790 202 3794
rect 204 3790 208 3794
rect 210 3790 214 3794
rect 216 3790 220 3794
rect 222 3790 226 3794
rect 228 3790 232 3794
rect 234 3790 238 3794
rect 240 3790 244 3794
rect 246 3790 250 3794
rect 252 3790 256 3794
rect 258 3790 262 3794
rect 264 3790 268 3794
rect 270 3790 274 3794
rect 276 3790 280 3794
rect 282 3790 286 3794
rect 288 3790 292 3794
rect 294 3790 298 3794
rect 300 3790 304 3794
rect 306 3790 310 3794
rect 312 3790 316 3794
rect 318 3790 322 3794
rect 324 3790 328 3794
rect 330 3790 334 3794
rect 336 3790 340 3794
rect 342 3790 346 3794
rect 348 3790 352 3794
rect 354 3790 358 3794
rect 360 3790 364 3794
rect 366 3790 370 3794
rect 372 3790 376 3794
rect 378 3790 382 3794
rect 384 3790 388 3794
rect 390 3790 394 3794
rect 396 3790 400 3794
rect 402 3790 406 3794
rect 408 3790 412 3794
rect 414 3790 418 3794
rect 420 3790 424 3794
rect 426 3790 430 3794
rect 432 3790 436 3794
rect 438 3790 442 3794
rect 444 3790 448 3794
rect 450 3790 454 3794
rect 456 3790 460 3794
rect 462 3790 466 3794
rect 468 3790 472 3794
rect 474 3790 478 3794
rect 480 3790 484 3794
rect 486 3790 490 3794
rect 492 3790 496 3794
rect 498 3790 502 3794
rect 504 3790 508 3794
rect 144 3784 148 3788
rect 144 3778 148 3782
rect 144 3772 148 3776
rect 144 3766 148 3770
rect 144 3760 148 3764
rect 144 3754 148 3758
rect 144 3748 148 3752
rect 144 3742 148 3746
rect 144 3736 148 3740
rect 144 3730 148 3734
rect 144 3724 148 3728
rect 144 3718 148 3722
rect 144 3712 148 3716
rect 144 3706 148 3710
rect 144 3700 148 3704
rect 144 3694 148 3698
rect 144 3688 148 3692
rect 144 3682 148 3686
rect 144 3676 148 3680
rect 144 3670 148 3674
rect 144 3664 148 3668
rect 144 3658 148 3662
rect 144 3652 148 3656
rect 144 3646 148 3650
rect 144 3640 148 3644
rect 144 3634 148 3638
rect 144 3628 148 3632
rect 144 3622 148 3626
rect 144 3616 148 3620
rect 144 3610 148 3614
rect 144 3604 148 3608
rect 144 3598 148 3602
rect 144 3592 148 3596
rect 144 3586 148 3590
rect 144 3580 148 3584
rect 144 3574 148 3578
rect 144 3568 148 3572
rect 144 3538 148 3542
rect 144 3532 148 3536
rect 144 3526 148 3530
rect 144 3520 148 3524
rect 144 3514 148 3518
rect 144 3508 148 3512
rect 144 3502 148 3506
rect 144 3496 148 3500
rect 144 3490 148 3494
rect 144 3484 148 3488
rect 144 3478 148 3482
rect 144 3472 148 3476
rect 144 3466 148 3470
rect 144 3460 148 3464
rect 144 3454 148 3458
rect 144 3448 148 3452
rect 144 3442 148 3446
rect 144 3436 148 3440
rect 144 3430 148 3434
rect 144 3424 148 3428
rect 144 3418 148 3422
rect 144 3412 148 3416
rect 144 3406 148 3410
rect 144 3400 148 3404
rect 144 3394 148 3398
rect 144 3388 148 3392
rect 144 3382 148 3386
rect 144 3376 148 3380
rect 144 3370 148 3374
rect 144 3364 148 3368
rect 144 3358 148 3362
rect 144 3352 148 3356
rect 144 3346 148 3350
rect 144 3340 148 3344
rect 144 3334 148 3338
rect 144 3328 148 3332
rect 144 3322 148 3326
rect 144 3316 148 3320
rect 150 3316 154 3320
rect 156 3316 160 3320
rect 162 3316 166 3320
rect 168 3316 172 3320
rect 174 3316 178 3320
rect 180 3316 184 3320
rect 186 3316 190 3320
rect 192 3316 196 3320
rect 198 3316 202 3320
rect 204 3316 208 3320
rect 210 3316 214 3320
rect 216 3316 220 3320
rect 222 3316 226 3320
rect 228 3316 232 3320
rect 234 3316 238 3320
rect 240 3316 244 3320
rect 246 3316 250 3320
rect 252 3316 256 3320
rect 258 3316 262 3320
rect 264 3316 268 3320
rect 270 3316 274 3320
rect 276 3316 280 3320
rect 282 3316 286 3320
rect 288 3316 292 3320
rect 294 3316 298 3320
rect 300 3316 304 3320
rect 306 3316 310 3320
rect 312 3316 316 3320
rect 318 3316 322 3320
rect 324 3316 328 3320
rect 330 3316 334 3320
rect 336 3316 340 3320
rect 342 3316 346 3320
rect 348 3316 352 3320
rect 354 3316 358 3320
rect 360 3316 364 3320
rect 366 3316 370 3320
rect 372 3316 376 3320
rect 378 3316 382 3320
rect 384 3316 388 3320
rect 390 3316 394 3320
rect 396 3316 400 3320
rect 402 3316 406 3320
rect 408 3316 412 3320
rect 414 3316 418 3320
rect 420 3316 424 3320
rect 426 3316 430 3320
rect 432 3316 436 3320
rect 438 3316 442 3320
rect 444 3316 448 3320
rect 450 3316 454 3320
rect 456 3316 460 3320
rect 462 3316 466 3320
rect 468 3316 472 3320
rect 474 3316 478 3320
rect 480 3316 484 3320
rect 486 3316 490 3320
rect 492 3316 496 3320
rect 498 3316 502 3320
rect 504 3316 508 3320
rect 144 3310 148 3314
rect 144 3304 148 3308
rect 144 3298 148 3302
rect 144 3292 148 3296
rect 144 3286 148 3290
rect 144 3280 148 3284
rect 144 3274 148 3278
rect 144 3268 148 3272
rect 144 3262 148 3266
rect 144 3256 148 3260
rect 144 3250 148 3254
rect 144 3244 148 3248
rect 144 3238 148 3242
rect 144 3232 148 3236
rect 144 3226 148 3230
rect 144 3220 148 3224
rect 144 3214 148 3218
rect 144 3208 148 3212
rect 144 3202 148 3206
rect 144 3196 148 3200
rect 144 3190 148 3194
rect 144 3184 148 3188
rect 144 3178 148 3182
rect 144 3172 148 3176
rect 144 3166 148 3170
rect 144 3160 148 3164
rect 144 3154 148 3158
rect 144 3148 148 3152
rect 144 3142 148 3146
rect 144 3136 148 3140
rect 144 3130 148 3134
rect 144 3124 148 3128
rect 144 3118 148 3122
rect 144 3112 148 3116
rect 144 3106 148 3110
rect 144 3100 148 3104
rect 144 3094 148 3098
rect 144 3064 148 3068
rect 144 3058 148 3062
rect 144 3052 148 3056
rect 144 3046 148 3050
rect 144 3040 148 3044
rect 144 3034 148 3038
rect 144 3028 148 3032
rect 144 3022 148 3026
rect 144 3016 148 3020
rect 144 3010 148 3014
rect 144 3004 148 3008
rect 144 2998 148 3002
rect 144 2992 148 2996
rect 144 2986 148 2990
rect 144 2980 148 2984
rect 144 2974 148 2978
rect 144 2968 148 2972
rect 144 2962 148 2966
rect 144 2956 148 2960
rect 144 2950 148 2954
rect 144 2944 148 2948
rect 144 2938 148 2942
rect 144 2932 148 2936
rect 144 2926 148 2930
rect 144 2920 148 2924
rect 144 2914 148 2918
rect 144 2908 148 2912
rect 144 2902 148 2906
rect 144 2896 148 2900
rect 144 2890 148 2894
rect 144 2884 148 2888
rect 144 2878 148 2882
rect 144 2872 148 2876
rect 144 2866 148 2870
rect 144 2860 148 2864
rect 144 2854 148 2858
rect 144 2848 148 2852
rect 144 2842 148 2846
rect 150 2842 154 2846
rect 156 2842 160 2846
rect 162 2842 166 2846
rect 168 2842 172 2846
rect 174 2842 178 2846
rect 180 2842 184 2846
rect 186 2842 190 2846
rect 192 2842 196 2846
rect 198 2842 202 2846
rect 204 2842 208 2846
rect 210 2842 214 2846
rect 216 2842 220 2846
rect 222 2842 226 2846
rect 228 2842 232 2846
rect 234 2842 238 2846
rect 240 2842 244 2846
rect 246 2842 250 2846
rect 252 2842 256 2846
rect 258 2842 262 2846
rect 264 2842 268 2846
rect 270 2842 274 2846
rect 276 2842 280 2846
rect 282 2842 286 2846
rect 288 2842 292 2846
rect 294 2842 298 2846
rect 300 2842 304 2846
rect 306 2842 310 2846
rect 312 2842 316 2846
rect 318 2842 322 2846
rect 324 2842 328 2846
rect 330 2842 334 2846
rect 336 2842 340 2846
rect 342 2842 346 2846
rect 348 2842 352 2846
rect 354 2842 358 2846
rect 360 2842 364 2846
rect 366 2842 370 2846
rect 372 2842 376 2846
rect 378 2842 382 2846
rect 384 2842 388 2846
rect 390 2842 394 2846
rect 396 2842 400 2846
rect 402 2842 406 2846
rect 408 2842 412 2846
rect 414 2842 418 2846
rect 420 2842 424 2846
rect 426 2842 430 2846
rect 432 2842 436 2846
rect 438 2842 442 2846
rect 444 2842 448 2846
rect 450 2842 454 2846
rect 456 2842 460 2846
rect 462 2842 466 2846
rect 468 2842 472 2846
rect 474 2842 478 2846
rect 480 2842 484 2846
rect 486 2842 490 2846
rect 492 2842 496 2846
rect 498 2842 502 2846
rect 504 2842 508 2846
rect 144 2836 148 2840
rect 144 2830 148 2834
rect 144 2824 148 2828
rect 144 2818 148 2822
rect 144 2812 148 2816
rect 144 2806 148 2810
rect 144 2800 148 2804
rect 144 2794 148 2798
rect 144 2788 148 2792
rect 144 2782 148 2786
rect 144 2776 148 2780
rect 144 2770 148 2774
rect 144 2764 148 2768
rect 144 2758 148 2762
rect 144 2752 148 2756
rect 144 2746 148 2750
rect 144 2740 148 2744
rect 144 2734 148 2738
rect 144 2728 148 2732
rect 144 2722 148 2726
rect 144 2716 148 2720
rect 144 2710 148 2714
rect 144 2704 148 2708
rect 144 2698 148 2702
rect 144 2692 148 2696
rect 144 2686 148 2690
rect 144 2680 148 2684
rect 144 2674 148 2678
rect 144 2668 148 2672
rect 144 2662 148 2666
rect 144 2656 148 2660
rect 144 2650 148 2654
rect 144 2644 148 2648
rect 144 2638 148 2642
rect 144 2632 148 2636
rect 144 2626 148 2630
rect 144 2620 148 2624
rect 144 2590 148 2594
rect 144 2584 148 2588
rect 144 2578 148 2582
rect 144 2572 148 2576
rect 144 2566 148 2570
rect 144 2560 148 2564
rect 144 2554 148 2558
rect 144 2548 148 2552
rect 144 2542 148 2546
rect 144 2536 148 2540
rect 144 2530 148 2534
rect 144 2524 148 2528
rect 144 2518 148 2522
rect 144 2512 148 2516
rect 144 2506 148 2510
rect 144 2500 148 2504
rect 144 2494 148 2498
rect 144 2488 148 2492
rect 144 2482 148 2486
rect 144 2476 148 2480
rect 144 2470 148 2474
rect 144 2464 148 2468
rect 144 2458 148 2462
rect 144 2452 148 2456
rect 144 2446 148 2450
rect 144 2440 148 2444
rect 144 2434 148 2438
rect 144 2428 148 2432
rect 144 2422 148 2426
rect 144 2416 148 2420
rect 144 2410 148 2414
rect 144 2404 148 2408
rect 144 2398 148 2402
rect 144 2392 148 2396
rect 144 2386 148 2390
rect 144 2380 148 2384
rect 144 2374 148 2378
rect 144 2368 148 2372
rect 150 2368 154 2372
rect 156 2368 160 2372
rect 162 2368 166 2372
rect 168 2368 172 2372
rect 174 2368 178 2372
rect 180 2368 184 2372
rect 186 2368 190 2372
rect 192 2368 196 2372
rect 198 2368 202 2372
rect 204 2368 208 2372
rect 210 2368 214 2372
rect 216 2368 220 2372
rect 222 2368 226 2372
rect 228 2368 232 2372
rect 234 2368 238 2372
rect 240 2368 244 2372
rect 246 2368 250 2372
rect 252 2368 256 2372
rect 258 2368 262 2372
rect 264 2368 268 2372
rect 270 2368 274 2372
rect 276 2368 280 2372
rect 282 2368 286 2372
rect 288 2368 292 2372
rect 294 2368 298 2372
rect 300 2368 304 2372
rect 306 2368 310 2372
rect 312 2368 316 2372
rect 318 2368 322 2372
rect 324 2368 328 2372
rect 330 2368 334 2372
rect 336 2368 340 2372
rect 342 2368 346 2372
rect 348 2368 352 2372
rect 354 2368 358 2372
rect 360 2368 364 2372
rect 366 2368 370 2372
rect 372 2368 376 2372
rect 378 2368 382 2372
rect 384 2368 388 2372
rect 390 2368 394 2372
rect 396 2368 400 2372
rect 402 2368 406 2372
rect 408 2368 412 2372
rect 414 2368 418 2372
rect 420 2368 424 2372
rect 426 2368 430 2372
rect 432 2368 436 2372
rect 438 2368 442 2372
rect 444 2368 448 2372
rect 450 2368 454 2372
rect 456 2368 460 2372
rect 462 2368 466 2372
rect 468 2368 472 2372
rect 474 2368 478 2372
rect 480 2368 484 2372
rect 486 2368 490 2372
rect 492 2368 496 2372
rect 498 2368 502 2372
rect 504 2368 508 2372
rect 144 2362 148 2366
rect 144 2356 148 2360
rect 144 2350 148 2354
rect 144 2344 148 2348
rect 144 2338 148 2342
rect 144 2332 148 2336
rect 144 2326 148 2330
rect 144 2320 148 2324
rect 144 2314 148 2318
rect 144 2308 148 2312
rect 144 2302 148 2306
rect 144 2296 148 2300
rect 144 2290 148 2294
rect 144 2284 148 2288
rect 144 2278 148 2282
rect 144 2272 148 2276
rect 144 2266 148 2270
rect 144 2260 148 2264
rect 144 2254 148 2258
rect 144 2248 148 2252
rect 144 2242 148 2246
rect 144 2236 148 2240
rect 144 2230 148 2234
rect 144 2224 148 2228
rect 144 2218 148 2222
rect 144 2212 148 2216
rect 144 2206 148 2210
rect 144 2200 148 2204
rect 144 2194 148 2198
rect 144 2188 148 2192
rect 144 2182 148 2186
rect 144 2176 148 2180
rect 144 2170 148 2174
rect 144 2164 148 2168
rect 144 2158 148 2162
rect 144 2152 148 2156
rect 144 2146 148 2150
rect 144 2116 148 2120
rect 144 2110 148 2114
rect 144 2104 148 2108
rect 144 2098 148 2102
rect 144 2092 148 2096
rect 144 2086 148 2090
rect 144 2080 148 2084
rect 144 2074 148 2078
rect 144 2068 148 2072
rect 144 2062 148 2066
rect 144 2056 148 2060
rect 144 2050 148 2054
rect 144 2044 148 2048
rect 144 2038 148 2042
rect 144 2032 148 2036
rect 144 2026 148 2030
rect 144 2020 148 2024
rect 144 2014 148 2018
rect 144 2008 148 2012
rect 144 2002 148 2006
rect 144 1996 148 2000
rect 144 1990 148 1994
rect 144 1984 148 1988
rect 144 1978 148 1982
rect 144 1972 148 1976
rect 144 1966 148 1970
rect 144 1960 148 1964
rect 144 1954 148 1958
rect 144 1948 148 1952
rect 144 1942 148 1946
rect 144 1936 148 1940
rect 144 1930 148 1934
rect 144 1924 148 1928
rect 144 1918 148 1922
rect 144 1912 148 1916
rect 144 1906 148 1910
rect 144 1900 148 1904
rect 144 1894 148 1898
rect 150 1894 154 1898
rect 156 1894 160 1898
rect 162 1894 166 1898
rect 168 1894 172 1898
rect 174 1894 178 1898
rect 180 1894 184 1898
rect 186 1894 190 1898
rect 192 1894 196 1898
rect 198 1894 202 1898
rect 204 1894 208 1898
rect 210 1894 214 1898
rect 216 1894 220 1898
rect 222 1894 226 1898
rect 228 1894 232 1898
rect 234 1894 238 1898
rect 240 1894 244 1898
rect 246 1894 250 1898
rect 252 1894 256 1898
rect 258 1894 262 1898
rect 264 1894 268 1898
rect 270 1894 274 1898
rect 276 1894 280 1898
rect 282 1894 286 1898
rect 288 1894 292 1898
rect 294 1894 298 1898
rect 300 1894 304 1898
rect 306 1894 310 1898
rect 312 1894 316 1898
rect 318 1894 322 1898
rect 324 1894 328 1898
rect 330 1894 334 1898
rect 336 1894 340 1898
rect 342 1894 346 1898
rect 348 1894 352 1898
rect 354 1894 358 1898
rect 360 1894 364 1898
rect 366 1894 370 1898
rect 372 1894 376 1898
rect 378 1894 382 1898
rect 384 1894 388 1898
rect 390 1894 394 1898
rect 396 1894 400 1898
rect 402 1894 406 1898
rect 408 1894 412 1898
rect 414 1894 418 1898
rect 420 1894 424 1898
rect 426 1894 430 1898
rect 432 1894 436 1898
rect 438 1894 442 1898
rect 444 1894 448 1898
rect 450 1894 454 1898
rect 456 1894 460 1898
rect 462 1894 466 1898
rect 468 1894 472 1898
rect 474 1894 478 1898
rect 480 1894 484 1898
rect 486 1894 490 1898
rect 492 1894 496 1898
rect 498 1894 502 1898
rect 504 1894 508 1898
rect 144 1888 148 1892
rect 144 1882 148 1886
rect 144 1876 148 1880
rect 144 1870 148 1874
rect 144 1864 148 1868
rect 144 1858 148 1862
rect 144 1852 148 1856
rect 144 1846 148 1850
rect 144 1840 148 1844
rect 144 1834 148 1838
rect 144 1828 148 1832
rect 144 1822 148 1826
rect 144 1816 148 1820
rect 144 1810 148 1814
rect 144 1804 148 1808
rect 144 1798 148 1802
rect 144 1792 148 1796
rect 144 1786 148 1790
rect 144 1780 148 1784
rect 144 1774 148 1778
rect 144 1768 148 1772
rect 144 1762 148 1766
rect 144 1756 148 1760
rect 144 1750 148 1754
rect 144 1744 148 1748
rect 144 1738 148 1742
rect 144 1732 148 1736
rect 144 1726 148 1730
rect 144 1720 148 1724
rect 144 1714 148 1718
rect 144 1708 148 1712
rect 144 1702 148 1706
rect 144 1696 148 1700
rect 144 1690 148 1694
rect 144 1684 148 1688
rect 144 1678 148 1682
rect 144 1672 148 1676
rect 144 1642 148 1646
rect 144 1636 148 1640
rect 144 1630 148 1634
rect 144 1624 148 1628
rect 144 1618 148 1622
rect 144 1612 148 1616
rect 144 1606 148 1610
rect 144 1600 148 1604
rect 144 1594 148 1598
rect 144 1588 148 1592
rect 144 1582 148 1586
rect 144 1576 148 1580
rect 144 1570 148 1574
rect 144 1564 148 1568
rect 144 1558 148 1562
rect 144 1552 148 1556
rect 144 1546 148 1550
rect 144 1540 148 1544
rect 144 1534 148 1538
rect 144 1528 148 1532
rect 144 1522 148 1526
rect 144 1516 148 1520
rect 144 1510 148 1514
rect 144 1504 148 1508
rect 144 1498 148 1502
rect 144 1492 148 1496
rect 144 1486 148 1490
rect 144 1480 148 1484
rect 144 1474 148 1478
rect 144 1468 148 1472
rect 144 1462 148 1466
rect 144 1456 148 1460
rect 144 1450 148 1454
rect 144 1444 148 1448
rect 144 1438 148 1442
rect 144 1432 148 1436
rect 144 1426 148 1430
rect 144 1420 148 1424
rect 150 1420 154 1424
rect 156 1420 160 1424
rect 162 1420 166 1424
rect 168 1420 172 1424
rect 174 1420 178 1424
rect 180 1420 184 1424
rect 186 1420 190 1424
rect 192 1420 196 1424
rect 198 1420 202 1424
rect 204 1420 208 1424
rect 210 1420 214 1424
rect 216 1420 220 1424
rect 222 1420 226 1424
rect 228 1420 232 1424
rect 234 1420 238 1424
rect 240 1420 244 1424
rect 246 1420 250 1424
rect 252 1420 256 1424
rect 258 1420 262 1424
rect 264 1420 268 1424
rect 270 1420 274 1424
rect 276 1420 280 1424
rect 282 1420 286 1424
rect 288 1420 292 1424
rect 294 1420 298 1424
rect 300 1420 304 1424
rect 306 1420 310 1424
rect 312 1420 316 1424
rect 318 1420 322 1424
rect 324 1420 328 1424
rect 330 1420 334 1424
rect 336 1420 340 1424
rect 342 1420 346 1424
rect 348 1420 352 1424
rect 354 1420 358 1424
rect 360 1420 364 1424
rect 366 1420 370 1424
rect 372 1420 376 1424
rect 378 1420 382 1424
rect 384 1420 388 1424
rect 390 1420 394 1424
rect 396 1420 400 1424
rect 402 1420 406 1424
rect 408 1420 412 1424
rect 414 1420 418 1424
rect 420 1420 424 1424
rect 426 1420 430 1424
rect 432 1420 436 1424
rect 438 1420 442 1424
rect 444 1420 448 1424
rect 450 1420 454 1424
rect 456 1420 460 1424
rect 462 1420 466 1424
rect 468 1420 472 1424
rect 474 1420 478 1424
rect 480 1420 484 1424
rect 486 1420 490 1424
rect 492 1420 496 1424
rect 498 1420 502 1424
rect 504 1420 508 1424
rect 144 1414 148 1418
rect 144 1408 148 1412
rect 144 1402 148 1406
rect 144 1396 148 1400
rect 144 1390 148 1394
rect 144 1384 148 1388
rect 144 1378 148 1382
rect 144 1372 148 1376
rect 144 1366 148 1370
rect 144 1360 148 1364
rect 144 1354 148 1358
rect 144 1348 148 1352
rect 144 1342 148 1346
rect 144 1336 148 1340
rect 144 1330 148 1334
rect 144 1324 148 1328
rect 144 1318 148 1322
rect 144 1312 148 1316
rect 144 1306 148 1310
rect 144 1300 148 1304
rect 144 1294 148 1298
rect 144 1288 148 1292
rect 144 1282 148 1286
rect 144 1276 148 1280
rect 144 1270 148 1274
rect 144 1264 148 1268
rect 144 1258 148 1262
rect 144 1252 148 1256
rect 144 1246 148 1250
rect 144 1240 148 1244
rect 144 1234 148 1238
rect 144 1228 148 1232
rect 144 1222 148 1226
rect 144 1216 148 1220
rect 144 1210 148 1214
rect 144 1204 148 1208
rect 144 1198 148 1202
rect 144 1168 148 1172
rect 144 1162 148 1166
rect 144 1156 148 1160
rect 144 1150 148 1154
rect 144 1144 148 1148
rect 144 1138 148 1142
rect 144 1132 148 1136
rect 144 1126 148 1130
rect 144 1120 148 1124
rect 144 1114 148 1118
rect 144 1108 148 1112
rect 144 1102 148 1106
rect 144 1096 148 1100
rect 144 1090 148 1094
rect 144 1084 148 1088
rect 144 1078 148 1082
rect 144 1072 148 1076
rect 144 1066 148 1070
rect 144 1060 148 1064
rect 144 1054 148 1058
rect 144 1048 148 1052
rect 144 1042 148 1046
rect 144 1036 148 1040
rect 144 1030 148 1034
rect 144 1024 148 1028
rect 144 1018 148 1022
rect 144 1012 148 1016
rect 144 1006 148 1010
rect 144 1000 148 1004
rect 144 994 148 998
rect 144 988 148 992
rect 144 982 148 986
rect 144 976 148 980
rect 144 970 148 974
rect 144 964 148 968
rect 144 958 148 962
rect 144 952 148 956
rect 144 946 148 950
rect 150 946 154 950
rect 156 946 160 950
rect 162 946 166 950
rect 168 946 172 950
rect 174 946 178 950
rect 180 946 184 950
rect 186 946 190 950
rect 192 946 196 950
rect 198 946 202 950
rect 204 946 208 950
rect 210 946 214 950
rect 216 946 220 950
rect 222 946 226 950
rect 228 946 232 950
rect 234 946 238 950
rect 240 946 244 950
rect 246 946 250 950
rect 252 946 256 950
rect 258 946 262 950
rect 264 946 268 950
rect 270 946 274 950
rect 276 946 280 950
rect 282 946 286 950
rect 288 946 292 950
rect 294 946 298 950
rect 300 946 304 950
rect 306 946 310 950
rect 312 946 316 950
rect 318 946 322 950
rect 324 946 328 950
rect 330 946 334 950
rect 336 946 340 950
rect 342 946 346 950
rect 348 946 352 950
rect 354 946 358 950
rect 360 946 364 950
rect 366 946 370 950
rect 372 946 376 950
rect 378 946 382 950
rect 384 946 388 950
rect 390 946 394 950
rect 396 946 400 950
rect 402 946 406 950
rect 408 946 412 950
rect 414 946 418 950
rect 420 946 424 950
rect 426 946 430 950
rect 432 946 436 950
rect 438 946 442 950
rect 444 946 448 950
rect 450 946 454 950
rect 456 946 460 950
rect 462 946 466 950
rect 468 946 472 950
rect 474 946 478 950
rect 480 946 484 950
rect 486 946 490 950
rect 492 946 496 950
rect 498 946 502 950
rect 504 946 508 950
rect 144 940 148 944
rect 144 934 148 938
rect 144 928 148 932
rect 144 922 148 926
rect 144 916 148 920
rect 144 910 148 914
rect 144 904 148 908
rect 144 898 148 902
rect 144 892 148 896
rect 144 886 148 890
rect 144 880 148 884
rect 144 874 148 878
rect 144 868 148 872
rect 144 862 148 866
rect 144 856 148 860
rect 144 850 148 854
rect 144 844 148 848
rect 144 838 148 842
rect 144 832 148 836
rect 144 826 148 830
rect 144 820 148 824
rect 144 814 148 818
rect 144 808 148 812
rect 144 802 148 806
rect 144 796 148 800
rect 144 790 148 794
rect 144 784 148 788
rect 144 778 148 782
rect 144 772 148 776
rect 144 766 148 770
rect 144 760 148 764
rect 144 754 148 758
rect 144 748 148 752
rect 144 742 148 746
rect 144 736 148 740
rect 144 730 148 734
rect 144 724 148 728
rect 144 694 148 698
rect 144 688 148 692
rect 144 682 148 686
rect 144 676 148 680
rect 144 670 148 674
rect 144 664 148 668
rect 144 658 148 662
rect 144 652 148 656
rect 144 646 148 650
rect 144 640 148 644
rect 144 634 148 638
rect 144 628 148 632
rect 144 622 148 626
rect 144 616 148 620
rect 144 610 148 614
rect 144 604 148 608
rect 144 598 148 602
rect 144 592 148 596
rect 144 586 148 590
rect 144 580 148 584
rect 144 574 148 578
rect 144 568 148 572
rect 144 562 148 566
rect 144 556 148 560
rect 144 550 148 554
rect 144 544 148 548
rect 144 538 148 542
rect 144 532 148 536
rect 144 526 148 530
rect 144 520 148 524
rect 144 514 148 518
rect 144 508 148 512
rect 144 502 148 506
rect 144 496 148 500
rect 144 490 148 494
rect 144 484 148 488
rect 144 478 148 482
rect 144 472 148 476
rect 150 472 154 476
rect 156 472 160 476
rect 162 472 166 476
rect 168 472 172 476
rect 174 472 178 476
rect 180 472 184 476
rect 186 472 190 476
rect 192 472 196 476
rect 198 472 202 476
rect 204 472 208 476
rect 210 472 214 476
rect 216 472 220 476
rect 222 472 226 476
rect 228 472 232 476
rect 234 472 238 476
rect 240 472 244 476
rect 246 472 250 476
rect 252 472 256 476
rect 258 472 262 476
rect 264 472 268 476
rect 270 472 274 476
rect 276 472 280 476
rect 282 472 286 476
rect 288 472 292 476
rect 294 472 298 476
rect 300 472 304 476
rect 306 472 310 476
rect 312 472 316 476
rect 318 472 322 476
rect 324 472 328 476
rect 330 472 334 476
rect 336 472 340 476
rect 342 472 346 476
rect 348 472 352 476
rect 354 472 358 476
rect 360 472 364 476
rect 366 472 370 476
rect 372 472 376 476
rect 378 472 382 476
rect 384 472 388 476
rect 390 472 394 476
rect 396 472 400 476
rect 402 472 406 476
rect 408 472 412 476
rect 414 472 418 476
rect 420 472 424 476
rect 426 472 430 476
rect 432 472 436 476
rect 438 472 442 476
rect 444 472 448 476
rect 450 472 454 476
rect 456 472 460 476
rect 462 472 466 476
rect 468 472 472 476
rect 474 472 478 476
rect 480 472 484 476
rect 486 472 490 476
rect 492 472 496 476
rect 498 472 502 476
rect 504 472 508 476
rect 144 466 148 470
rect 144 460 148 464
rect 144 454 148 458
rect 144 448 148 452
rect 144 442 148 446
rect 144 436 148 440
rect 144 430 148 434
rect 144 424 148 428
rect 144 418 148 422
rect 144 412 148 416
rect 144 406 148 410
rect 144 400 148 404
rect 144 394 148 398
rect 144 388 148 392
rect 144 382 148 386
rect 144 376 148 380
rect 144 370 148 374
rect 144 364 148 368
rect 144 358 148 362
rect 144 352 148 356
rect 144 346 148 350
rect 144 340 148 344
rect 144 334 148 338
rect 144 328 148 332
rect 144 322 148 326
rect 144 316 148 320
rect 144 310 148 314
rect 144 304 148 308
rect 144 298 148 302
rect 144 292 148 296
rect 144 286 148 290
rect 144 280 148 284
rect 144 274 148 278
rect 144 268 148 272
rect 144 262 148 266
rect 144 256 148 260
rect 144 250 148 254
rect 144 220 148 224
rect 144 214 148 218
rect 144 208 148 212
rect 144 202 148 206
rect 144 196 148 200
rect 144 190 148 194
rect 144 184 148 188
rect 144 178 148 182
rect 144 172 148 176
rect 144 166 148 170
rect 144 160 148 164
rect 144 154 148 158
rect 144 148 148 152
rect 144 142 148 146
rect 144 136 148 140
rect 144 130 148 134
rect 144 124 148 128
rect 144 118 148 122
rect 144 112 148 116
rect 144 106 148 110
rect 144 100 148 104
rect 144 94 148 98
rect 144 88 148 92
rect 144 82 148 86
rect 144 76 148 80
rect 144 70 148 74
rect 144 64 148 68
rect 144 58 148 62
rect 144 52 148 56
rect 144 46 148 50
rect 144 40 148 44
rect 144 34 148 38
rect 144 28 148 32
rect 144 22 148 26
rect 144 16 148 20
rect 144 10 148 14
rect 144 4 148 8
<< polysilicon >>
rect 7 4138 142 4262
rect 7 4134 137 4138
rect 141 4134 142 4138
rect 7 4132 142 4134
rect 7 4128 137 4132
rect 141 4128 142 4132
rect 7 4126 142 4128
rect 7 4122 137 4126
rect 141 4122 142 4126
rect 7 4120 142 4122
rect 7 4116 137 4120
rect 141 4116 142 4120
rect 7 4114 142 4116
rect 7 4110 137 4114
rect 141 4110 142 4114
rect 7 4108 142 4110
rect 7 4104 137 4108
rect 141 4104 142 4108
rect 7 4102 142 4104
rect 7 4098 137 4102
rect 141 4098 142 4102
rect 7 3960 142 4098
rect 7 3956 8 3960
rect 12 3956 137 3960
rect 141 3956 142 3960
rect 7 3954 142 3956
rect 7 3950 8 3954
rect 12 3950 137 3954
rect 141 3950 142 3954
rect 7 3948 142 3950
rect 7 3944 8 3948
rect 12 3944 137 3948
rect 141 3944 142 3948
rect 7 3942 142 3944
rect 7 3938 8 3942
rect 12 3938 137 3942
rect 141 3938 142 3942
rect 7 3936 142 3938
rect 7 3932 8 3936
rect 12 3932 137 3936
rect 141 3932 142 3936
rect 7 3930 142 3932
rect 7 3926 8 3930
rect 12 3926 137 3930
rect 141 3926 142 3930
rect 7 3924 142 3926
rect 7 3920 8 3924
rect 12 3920 137 3924
rect 141 3920 142 3924
rect 7 3664 142 3920
rect 7 3660 8 3664
rect 12 3660 137 3664
rect 141 3660 142 3664
rect 7 3658 142 3660
rect 7 3654 8 3658
rect 12 3654 137 3658
rect 141 3654 142 3658
rect 7 3652 142 3654
rect 7 3648 8 3652
rect 12 3648 137 3652
rect 141 3648 142 3652
rect 7 3646 142 3648
rect 7 3642 8 3646
rect 12 3642 137 3646
rect 141 3642 142 3646
rect 7 3640 142 3642
rect 7 3636 8 3640
rect 12 3636 137 3640
rect 141 3636 142 3640
rect 7 3634 142 3636
rect 7 3630 8 3634
rect 12 3630 137 3634
rect 141 3630 142 3634
rect 7 3628 142 3630
rect 7 3624 8 3628
rect 12 3624 137 3628
rect 141 3624 142 3628
rect 7 3486 142 3624
rect 7 3482 8 3486
rect 12 3482 137 3486
rect 141 3482 142 3486
rect 7 3480 142 3482
rect 7 3476 8 3480
rect 12 3476 137 3480
rect 141 3476 142 3480
rect 7 3474 142 3476
rect 7 3470 8 3474
rect 12 3470 137 3474
rect 141 3470 142 3474
rect 7 3468 142 3470
rect 7 3464 8 3468
rect 12 3464 137 3468
rect 141 3464 142 3468
rect 7 3462 142 3464
rect 7 3458 8 3462
rect 12 3458 137 3462
rect 141 3458 142 3462
rect 7 3456 142 3458
rect 7 3452 8 3456
rect 12 3452 137 3456
rect 141 3452 142 3456
rect 7 3450 142 3452
rect 7 3446 8 3450
rect 12 3446 137 3450
rect 141 3446 142 3450
rect 7 3190 142 3446
rect 7 3186 8 3190
rect 12 3186 137 3190
rect 141 3186 142 3190
rect 7 3184 142 3186
rect 7 3180 8 3184
rect 12 3180 137 3184
rect 141 3180 142 3184
rect 7 3178 142 3180
rect 7 3174 8 3178
rect 12 3174 137 3178
rect 141 3174 142 3178
rect 7 3172 142 3174
rect 7 3168 8 3172
rect 12 3168 137 3172
rect 141 3168 142 3172
rect 7 3166 142 3168
rect 7 3162 8 3166
rect 12 3162 137 3166
rect 141 3162 142 3166
rect 7 3160 142 3162
rect 7 3156 8 3160
rect 12 3156 137 3160
rect 141 3156 142 3160
rect 7 3154 142 3156
rect 7 3150 8 3154
rect 12 3150 137 3154
rect 141 3150 142 3154
rect 7 3012 142 3150
rect 7 3008 8 3012
rect 12 3008 137 3012
rect 141 3008 142 3012
rect 7 3006 142 3008
rect 7 3002 8 3006
rect 12 3002 137 3006
rect 141 3002 142 3006
rect 7 3000 142 3002
rect 7 2996 8 3000
rect 12 2996 137 3000
rect 141 2996 142 3000
rect 7 2994 142 2996
rect 7 2990 8 2994
rect 12 2990 137 2994
rect 141 2990 142 2994
rect 7 2988 142 2990
rect 7 2984 8 2988
rect 12 2984 137 2988
rect 141 2984 142 2988
rect 7 2982 142 2984
rect 7 2978 8 2982
rect 12 2978 137 2982
rect 141 2978 142 2982
rect 7 2976 142 2978
rect 7 2972 8 2976
rect 12 2972 137 2976
rect 141 2972 142 2976
rect 7 2716 142 2972
rect 7 2712 8 2716
rect 12 2712 137 2716
rect 141 2712 142 2716
rect 7 2710 142 2712
rect 7 2706 8 2710
rect 12 2706 137 2710
rect 141 2706 142 2710
rect 7 2704 142 2706
rect 7 2700 8 2704
rect 12 2700 137 2704
rect 141 2700 142 2704
rect 7 2698 142 2700
rect 7 2694 8 2698
rect 12 2694 137 2698
rect 141 2694 142 2698
rect 7 2692 142 2694
rect 7 2688 8 2692
rect 12 2688 137 2692
rect 141 2688 142 2692
rect 7 2686 142 2688
rect 7 2682 8 2686
rect 12 2682 137 2686
rect 141 2682 142 2686
rect 7 2680 142 2682
rect 7 2676 8 2680
rect 12 2676 137 2680
rect 141 2676 142 2680
rect 7 2538 142 2676
rect 7 2534 8 2538
rect 12 2534 137 2538
rect 141 2534 142 2538
rect 7 2532 142 2534
rect 7 2528 8 2532
rect 12 2528 137 2532
rect 141 2528 142 2532
rect 7 2526 142 2528
rect 7 2522 8 2526
rect 12 2522 137 2526
rect 141 2522 142 2526
rect 7 2520 142 2522
rect 7 2516 8 2520
rect 12 2516 137 2520
rect 141 2516 142 2520
rect 7 2514 142 2516
rect 7 2510 8 2514
rect 12 2510 137 2514
rect 141 2510 142 2514
rect 7 2508 142 2510
rect 7 2504 8 2508
rect 12 2504 137 2508
rect 141 2504 142 2508
rect 7 2502 142 2504
rect 7 2498 8 2502
rect 12 2498 137 2502
rect 141 2498 142 2502
rect 7 2242 142 2498
rect 7 2238 8 2242
rect 12 2238 137 2242
rect 141 2238 142 2242
rect 7 2236 142 2238
rect 7 2232 8 2236
rect 12 2232 137 2236
rect 141 2232 142 2236
rect 7 2230 142 2232
rect 7 2226 8 2230
rect 12 2226 137 2230
rect 141 2226 142 2230
rect 7 2224 142 2226
rect 7 2220 8 2224
rect 12 2220 137 2224
rect 141 2220 142 2224
rect 7 2218 142 2220
rect 7 2214 8 2218
rect 12 2214 137 2218
rect 141 2214 142 2218
rect 7 2212 142 2214
rect 7 2208 8 2212
rect 12 2208 137 2212
rect 141 2208 142 2212
rect 7 2206 142 2208
rect 7 2202 8 2206
rect 12 2202 137 2206
rect 141 2202 142 2206
rect 7 2064 142 2202
rect 7 2060 8 2064
rect 12 2060 137 2064
rect 141 2060 142 2064
rect 7 2058 142 2060
rect 7 2054 8 2058
rect 12 2054 137 2058
rect 141 2054 142 2058
rect 7 2052 142 2054
rect 7 2048 8 2052
rect 12 2048 137 2052
rect 141 2048 142 2052
rect 7 2046 142 2048
rect 7 2042 8 2046
rect 12 2042 137 2046
rect 141 2042 142 2046
rect 7 2040 142 2042
rect 7 2036 8 2040
rect 12 2036 137 2040
rect 141 2036 142 2040
rect 7 2034 142 2036
rect 7 2030 8 2034
rect 12 2030 137 2034
rect 141 2030 142 2034
rect 7 2028 142 2030
rect 7 2024 8 2028
rect 12 2024 137 2028
rect 141 2024 142 2028
rect 7 1768 142 2024
rect 7 1764 8 1768
rect 12 1764 137 1768
rect 141 1764 142 1768
rect 7 1762 142 1764
rect 7 1758 8 1762
rect 12 1758 137 1762
rect 141 1758 142 1762
rect 7 1756 142 1758
rect 7 1752 8 1756
rect 12 1752 137 1756
rect 141 1752 142 1756
rect 7 1750 142 1752
rect 7 1746 8 1750
rect 12 1746 137 1750
rect 141 1746 142 1750
rect 7 1744 142 1746
rect 7 1740 8 1744
rect 12 1740 137 1744
rect 141 1740 142 1744
rect 7 1738 142 1740
rect 7 1734 8 1738
rect 12 1734 137 1738
rect 141 1734 142 1738
rect 7 1732 142 1734
rect 7 1728 8 1732
rect 12 1728 137 1732
rect 141 1728 142 1732
rect 7 1590 142 1728
rect 7 1586 8 1590
rect 12 1586 137 1590
rect 141 1586 142 1590
rect 7 1584 142 1586
rect 7 1580 8 1584
rect 12 1580 137 1584
rect 141 1580 142 1584
rect 7 1578 142 1580
rect 7 1574 8 1578
rect 12 1574 137 1578
rect 141 1574 142 1578
rect 7 1572 142 1574
rect 7 1568 8 1572
rect 12 1568 137 1572
rect 141 1568 142 1572
rect 7 1566 142 1568
rect 7 1562 8 1566
rect 12 1562 137 1566
rect 141 1562 142 1566
rect 7 1560 142 1562
rect 7 1556 8 1560
rect 12 1556 137 1560
rect 141 1556 142 1560
rect 7 1554 142 1556
rect 7 1550 8 1554
rect 12 1550 137 1554
rect 141 1550 142 1554
rect 7 1294 142 1550
rect 7 1290 8 1294
rect 12 1290 137 1294
rect 141 1290 142 1294
rect 7 1288 142 1290
rect 7 1284 8 1288
rect 12 1284 137 1288
rect 141 1284 142 1288
rect 7 1282 142 1284
rect 7 1278 8 1282
rect 12 1278 137 1282
rect 141 1278 142 1282
rect 7 1276 142 1278
rect 7 1272 8 1276
rect 12 1272 137 1276
rect 141 1272 142 1276
rect 7 1270 142 1272
rect 7 1266 8 1270
rect 12 1266 137 1270
rect 141 1266 142 1270
rect 7 1264 142 1266
rect 7 1260 8 1264
rect 12 1260 137 1264
rect 141 1260 142 1264
rect 7 1258 142 1260
rect 7 1254 8 1258
rect 12 1254 137 1258
rect 141 1254 142 1258
rect 7 1116 142 1254
rect 7 1112 8 1116
rect 12 1112 137 1116
rect 141 1112 142 1116
rect 7 1110 142 1112
rect 7 1106 8 1110
rect 12 1106 137 1110
rect 141 1106 142 1110
rect 7 1104 142 1106
rect 7 1100 8 1104
rect 12 1100 137 1104
rect 141 1100 142 1104
rect 7 1098 142 1100
rect 7 1094 8 1098
rect 12 1094 137 1098
rect 141 1094 142 1098
rect 7 1092 142 1094
rect 7 1088 8 1092
rect 12 1088 137 1092
rect 141 1088 142 1092
rect 7 1086 142 1088
rect 7 1082 8 1086
rect 12 1082 137 1086
rect 141 1082 142 1086
rect 7 1080 142 1082
rect 7 1076 8 1080
rect 12 1076 137 1080
rect 141 1076 142 1080
rect 7 820 142 1076
rect 7 816 8 820
rect 12 816 137 820
rect 141 816 142 820
rect 7 814 142 816
rect 7 810 8 814
rect 12 810 137 814
rect 141 810 142 814
rect 7 808 142 810
rect 7 804 8 808
rect 12 804 137 808
rect 141 804 142 808
rect 7 802 142 804
rect 7 798 8 802
rect 12 798 137 802
rect 141 798 142 802
rect 7 796 142 798
rect 7 792 8 796
rect 12 792 137 796
rect 141 792 142 796
rect 7 790 142 792
rect 7 786 8 790
rect 12 786 137 790
rect 141 786 142 790
rect 7 784 142 786
rect 7 780 8 784
rect 12 780 137 784
rect 141 780 142 784
rect 7 642 142 780
rect 7 638 8 642
rect 12 638 137 642
rect 141 638 142 642
rect 7 636 142 638
rect 7 632 8 636
rect 12 632 137 636
rect 141 632 142 636
rect 7 630 142 632
rect 7 626 8 630
rect 12 626 137 630
rect 141 626 142 630
rect 7 624 142 626
rect 7 620 8 624
rect 12 620 137 624
rect 141 620 142 624
rect 7 618 142 620
rect 7 614 8 618
rect 12 614 137 618
rect 141 614 142 618
rect 7 612 142 614
rect 7 608 8 612
rect 12 608 137 612
rect 141 608 142 612
rect 7 606 142 608
rect 7 602 8 606
rect 12 602 137 606
rect 141 602 142 606
rect 7 346 142 602
rect 7 342 8 346
rect 12 342 137 346
rect 141 342 142 346
rect 7 340 142 342
rect 7 336 8 340
rect 12 336 137 340
rect 141 336 142 340
rect 7 334 142 336
rect 7 330 8 334
rect 12 330 137 334
rect 141 330 142 334
rect 7 328 142 330
rect 7 324 8 328
rect 12 324 137 328
rect 141 324 142 328
rect 7 322 142 324
rect 7 318 8 322
rect 12 318 137 322
rect 141 318 142 322
rect 7 316 142 318
rect 7 312 8 316
rect 12 312 137 316
rect 141 312 142 316
rect 7 310 142 312
rect 7 306 8 310
rect 12 306 137 310
rect 141 306 142 310
rect 7 168 142 306
rect 7 164 137 168
rect 141 164 142 168
rect 7 162 142 164
rect 7 158 137 162
rect 141 158 142 162
rect 7 156 142 158
rect 7 152 137 156
rect 141 152 142 156
rect 7 150 142 152
rect 7 146 137 150
rect 141 146 142 150
rect 7 144 142 146
rect 7 140 137 144
rect 141 140 142 144
rect 7 138 142 140
rect 7 134 137 138
rect 141 134 142 138
rect 7 132 142 134
rect 7 128 137 132
rect 141 128 142 132
rect 7 4 142 128
<< polycontact >>
rect 137 4134 141 4138
rect 137 4128 141 4132
rect 137 4122 141 4126
rect 137 4116 141 4120
rect 137 4110 141 4114
rect 137 4104 141 4108
rect 137 4098 141 4102
rect 8 3956 12 3960
rect 137 3956 141 3960
rect 8 3950 12 3954
rect 137 3950 141 3954
rect 8 3944 12 3948
rect 137 3944 141 3948
rect 8 3938 12 3942
rect 137 3938 141 3942
rect 8 3932 12 3936
rect 137 3932 141 3936
rect 8 3926 12 3930
rect 137 3926 141 3930
rect 8 3920 12 3924
rect 137 3920 141 3924
rect 8 3660 12 3664
rect 137 3660 141 3664
rect 8 3654 12 3658
rect 137 3654 141 3658
rect 8 3648 12 3652
rect 137 3648 141 3652
rect 8 3642 12 3646
rect 137 3642 141 3646
rect 8 3636 12 3640
rect 137 3636 141 3640
rect 8 3630 12 3634
rect 137 3630 141 3634
rect 8 3624 12 3628
rect 137 3624 141 3628
rect 8 3482 12 3486
rect 137 3482 141 3486
rect 8 3476 12 3480
rect 137 3476 141 3480
rect 8 3470 12 3474
rect 137 3470 141 3474
rect 8 3464 12 3468
rect 137 3464 141 3468
rect 8 3458 12 3462
rect 137 3458 141 3462
rect 8 3452 12 3456
rect 137 3452 141 3456
rect 8 3446 12 3450
rect 137 3446 141 3450
rect 8 3186 12 3190
rect 137 3186 141 3190
rect 8 3180 12 3184
rect 137 3180 141 3184
rect 8 3174 12 3178
rect 137 3174 141 3178
rect 8 3168 12 3172
rect 137 3168 141 3172
rect 8 3162 12 3166
rect 137 3162 141 3166
rect 8 3156 12 3160
rect 137 3156 141 3160
rect 8 3150 12 3154
rect 137 3150 141 3154
rect 8 3008 12 3012
rect 137 3008 141 3012
rect 8 3002 12 3006
rect 137 3002 141 3006
rect 8 2996 12 3000
rect 137 2996 141 3000
rect 8 2990 12 2994
rect 137 2990 141 2994
rect 8 2984 12 2988
rect 137 2984 141 2988
rect 8 2978 12 2982
rect 137 2978 141 2982
rect 8 2972 12 2976
rect 137 2972 141 2976
rect 8 2712 12 2716
rect 137 2712 141 2716
rect 8 2706 12 2710
rect 137 2706 141 2710
rect 8 2700 12 2704
rect 137 2700 141 2704
rect 8 2694 12 2698
rect 137 2694 141 2698
rect 8 2688 12 2692
rect 137 2688 141 2692
rect 8 2682 12 2686
rect 137 2682 141 2686
rect 8 2676 12 2680
rect 137 2676 141 2680
rect 8 2534 12 2538
rect 137 2534 141 2538
rect 8 2528 12 2532
rect 137 2528 141 2532
rect 8 2522 12 2526
rect 137 2522 141 2526
rect 8 2516 12 2520
rect 137 2516 141 2520
rect 8 2510 12 2514
rect 137 2510 141 2514
rect 8 2504 12 2508
rect 137 2504 141 2508
rect 8 2498 12 2502
rect 137 2498 141 2502
rect 8 2238 12 2242
rect 137 2238 141 2242
rect 8 2232 12 2236
rect 137 2232 141 2236
rect 8 2226 12 2230
rect 137 2226 141 2230
rect 8 2220 12 2224
rect 137 2220 141 2224
rect 8 2214 12 2218
rect 137 2214 141 2218
rect 8 2208 12 2212
rect 137 2208 141 2212
rect 8 2202 12 2206
rect 137 2202 141 2206
rect 8 2060 12 2064
rect 137 2060 141 2064
rect 8 2054 12 2058
rect 137 2054 141 2058
rect 8 2048 12 2052
rect 137 2048 141 2052
rect 8 2042 12 2046
rect 137 2042 141 2046
rect 8 2036 12 2040
rect 137 2036 141 2040
rect 8 2030 12 2034
rect 137 2030 141 2034
rect 8 2024 12 2028
rect 137 2024 141 2028
rect 8 1764 12 1768
rect 137 1764 141 1768
rect 8 1758 12 1762
rect 137 1758 141 1762
rect 8 1752 12 1756
rect 137 1752 141 1756
rect 8 1746 12 1750
rect 137 1746 141 1750
rect 8 1740 12 1744
rect 137 1740 141 1744
rect 8 1734 12 1738
rect 137 1734 141 1738
rect 8 1728 12 1732
rect 137 1728 141 1732
rect 8 1586 12 1590
rect 137 1586 141 1590
rect 8 1580 12 1584
rect 137 1580 141 1584
rect 8 1574 12 1578
rect 137 1574 141 1578
rect 8 1568 12 1572
rect 137 1568 141 1572
rect 8 1562 12 1566
rect 137 1562 141 1566
rect 8 1556 12 1560
rect 137 1556 141 1560
rect 8 1550 12 1554
rect 137 1550 141 1554
rect 8 1290 12 1294
rect 137 1290 141 1294
rect 8 1284 12 1288
rect 137 1284 141 1288
rect 8 1278 12 1282
rect 137 1278 141 1282
rect 8 1272 12 1276
rect 137 1272 141 1276
rect 8 1266 12 1270
rect 137 1266 141 1270
rect 8 1260 12 1264
rect 137 1260 141 1264
rect 8 1254 12 1258
rect 137 1254 141 1258
rect 8 1112 12 1116
rect 137 1112 141 1116
rect 8 1106 12 1110
rect 137 1106 141 1110
rect 8 1100 12 1104
rect 137 1100 141 1104
rect 8 1094 12 1098
rect 137 1094 141 1098
rect 8 1088 12 1092
rect 137 1088 141 1092
rect 8 1082 12 1086
rect 137 1082 141 1086
rect 8 1076 12 1080
rect 137 1076 141 1080
rect 8 816 12 820
rect 137 816 141 820
rect 8 810 12 814
rect 137 810 141 814
rect 8 804 12 808
rect 137 804 141 808
rect 8 798 12 802
rect 137 798 141 802
rect 8 792 12 796
rect 137 792 141 796
rect 8 786 12 790
rect 137 786 141 790
rect 8 780 12 784
rect 137 780 141 784
rect 8 638 12 642
rect 137 638 141 642
rect 8 632 12 636
rect 137 632 141 636
rect 8 626 12 630
rect 137 626 141 630
rect 8 620 12 624
rect 137 620 141 624
rect 8 614 12 618
rect 137 614 141 618
rect 8 608 12 612
rect 137 608 141 612
rect 8 602 12 606
rect 137 602 141 606
rect 8 342 12 346
rect 137 342 141 346
rect 8 336 12 340
rect 137 336 141 340
rect 8 330 12 334
rect 137 330 141 334
rect 8 324 12 328
rect 137 324 141 328
rect 8 318 12 322
rect 137 318 141 322
rect 8 312 12 316
rect 137 312 141 316
rect 8 306 12 310
rect 137 306 141 310
rect 137 164 141 168
rect 137 158 141 162
rect 137 152 141 156
rect 137 146 141 150
rect 137 140 141 144
rect 137 134 141 138
rect 137 128 141 132
<< metal1 >>
rect 144 4262 148 4264
rect 144 4256 148 4258
rect 144 4250 148 4252
rect 144 4244 148 4246
rect 144 4238 148 4240
rect 144 4232 148 4234
rect 144 4226 148 4228
rect 144 4220 148 4222
rect 144 4214 148 4216
rect 144 4208 148 4210
rect 144 4202 148 4204
rect 144 4196 148 4198
rect 144 4190 148 4192
rect 144 4184 148 4186
rect 144 4178 148 4180
rect 144 4172 148 4174
rect 144 4166 148 4168
rect 144 4160 148 4162
rect 144 4154 148 4156
rect 144 4148 148 4150
rect 144 4142 148 4144
rect 62 4134 63 4138
rect 72 4134 74 4138
rect 78 4134 80 4138
rect 84 4134 86 4138
rect 90 4134 92 4138
rect 101 4134 137 4138
rect 141 4136 148 4138
rect 141 4134 144 4136
rect 62 4132 144 4134
rect 62 4128 63 4132
rect 72 4128 74 4132
rect 78 4128 80 4132
rect 84 4128 86 4132
rect 90 4128 92 4132
rect 101 4128 137 4132
rect 141 4130 148 4132
rect 141 4128 144 4130
rect 62 4126 144 4128
rect 62 4122 63 4126
rect 72 4122 74 4126
rect 78 4122 80 4126
rect 84 4122 86 4126
rect 90 4122 92 4126
rect 101 4122 137 4126
rect 141 4124 148 4126
rect 141 4122 144 4124
rect 62 4120 144 4122
rect 62 4116 63 4120
rect 72 4116 74 4120
rect 78 4116 80 4120
rect 84 4116 86 4120
rect 90 4116 92 4120
rect 101 4116 137 4120
rect 141 4118 148 4120
rect 141 4116 144 4118
rect 62 4114 144 4116
rect 62 4110 63 4114
rect 72 4110 74 4114
rect 78 4110 80 4114
rect 84 4110 86 4114
rect 90 4110 92 4114
rect 101 4110 137 4114
rect 141 4112 148 4114
rect 141 4110 144 4112
rect 62 4108 144 4110
rect 62 4104 63 4108
rect 72 4104 74 4108
rect 78 4104 80 4108
rect 84 4104 86 4108
rect 90 4104 92 4108
rect 101 4104 137 4108
rect 141 4106 148 4108
rect 141 4104 144 4106
rect 62 4102 144 4104
rect 62 4098 63 4102
rect 72 4098 74 4102
rect 78 4098 80 4102
rect 84 4098 86 4102
rect 90 4098 92 4102
rect 101 4098 137 4102
rect 141 4100 148 4102
rect 141 4098 144 4100
rect 144 4094 148 4096
rect 4 4090 14 4094
rect 18 4090 20 4094
rect 24 4090 26 4094
rect 30 4090 32 4094
rect 36 4090 38 4094
rect 42 4090 43 4094
rect 47 4093 100 4094
rect 47 4090 64 4093
rect 0 4089 64 4090
rect 68 4089 70 4093
rect 74 4089 76 4093
rect 80 4089 82 4093
rect 86 4089 89 4093
rect 93 4089 95 4093
rect 99 4089 100 4093
rect 0 4088 100 4089
rect 4 4084 14 4088
rect 18 4084 20 4088
rect 24 4084 26 4088
rect 30 4084 32 4088
rect 36 4084 38 4088
rect 42 4084 43 4088
rect 47 4087 100 4088
rect 47 4084 64 4087
rect 0 4083 64 4084
rect 68 4083 70 4087
rect 74 4083 76 4087
rect 80 4083 82 4087
rect 86 4083 89 4087
rect 93 4083 95 4087
rect 99 4083 100 4087
rect 0 4082 100 4083
rect 4 4078 14 4082
rect 18 4078 20 4082
rect 24 4078 26 4082
rect 30 4078 32 4082
rect 36 4078 38 4082
rect 42 4078 43 4082
rect 47 4081 100 4082
rect 47 4078 64 4081
rect 0 4077 64 4078
rect 68 4077 70 4081
rect 74 4077 76 4081
rect 80 4077 82 4081
rect 86 4077 89 4081
rect 93 4077 95 4081
rect 99 4077 100 4081
rect 0 4076 100 4077
rect 4 4072 14 4076
rect 18 4072 20 4076
rect 24 4072 26 4076
rect 30 4072 32 4076
rect 36 4072 38 4076
rect 42 4072 43 4076
rect 47 4075 100 4076
rect 47 4072 64 4075
rect 0 4071 64 4072
rect 68 4071 70 4075
rect 74 4071 76 4075
rect 80 4071 82 4075
rect 86 4071 89 4075
rect 93 4071 95 4075
rect 99 4071 100 4075
rect 0 4070 100 4071
rect 4 4066 14 4070
rect 18 4066 20 4070
rect 24 4066 26 4070
rect 30 4066 32 4070
rect 36 4066 38 4070
rect 42 4066 43 4070
rect 47 4069 100 4070
rect 47 4066 64 4069
rect 0 4065 64 4066
rect 68 4065 70 4069
rect 74 4065 76 4069
rect 80 4065 82 4069
rect 86 4065 89 4069
rect 93 4065 95 4069
rect 99 4065 100 4069
rect 0 4064 100 4065
rect 111 4090 112 4094
rect 116 4090 119 4094
rect 123 4090 125 4094
rect 107 4088 129 4090
rect 144 4088 148 4090
rect 111 4084 112 4088
rect 116 4084 119 4088
rect 123 4084 125 4088
rect 129 4084 131 4088
rect 107 4082 135 4084
rect 111 4078 112 4082
rect 116 4078 119 4082
rect 123 4078 125 4082
rect 129 4078 131 4082
rect 107 4076 135 4078
rect 111 4072 112 4076
rect 116 4072 119 4076
rect 123 4072 125 4076
rect 129 4072 131 4076
rect 107 4070 135 4072
rect 111 4066 112 4070
rect 116 4066 119 4070
rect 123 4066 125 4070
rect 129 4066 131 4070
rect 107 4064 135 4066
rect 4 4060 14 4064
rect 18 4060 20 4064
rect 24 4060 26 4064
rect 30 4060 32 4064
rect 36 4060 38 4064
rect 42 4060 43 4064
rect 47 4060 48 4064
rect 111 4060 112 4064
rect 116 4060 119 4064
rect 123 4060 125 4064
rect 129 4060 131 4064
rect 0 4058 48 4060
rect 4 4054 14 4058
rect 18 4054 20 4058
rect 24 4054 26 4058
rect 30 4054 32 4058
rect 36 4054 38 4058
rect 42 4054 43 4058
rect 47 4054 48 4058
rect 52 4056 53 4060
rect 57 4056 58 4060
rect 52 4055 58 4056
rect 52 4051 53 4055
rect 57 4051 58 4055
rect 107 4058 135 4060
rect 111 4054 112 4058
rect 116 4054 119 4058
rect 123 4054 125 4058
rect 129 4054 131 4058
rect 144 4082 148 4084
rect 144 4076 148 4078
rect 144 4070 148 4072
rect 144 4064 148 4066
rect 144 4058 148 4060
rect 52 4050 58 4051
rect 4 4046 53 4050
rect 57 4046 58 4050
rect 4 4045 58 4046
rect 4 4041 53 4045
rect 57 4041 58 4045
rect 144 4052 148 4054
rect 144 4046 148 4048
rect 4 4013 53 4017
rect 57 4013 58 4017
rect 4 4012 58 4013
rect 4 4008 53 4012
rect 57 4008 58 4012
rect 52 4007 58 4008
rect 4 4000 14 4004
rect 18 4000 20 4004
rect 24 4000 26 4004
rect 30 4000 32 4004
rect 36 4000 38 4004
rect 42 4000 43 4004
rect 47 4000 48 4004
rect 0 3998 48 4000
rect 52 4003 53 4007
rect 57 4003 58 4007
rect 144 4010 148 4012
rect 144 4004 148 4006
rect 52 4002 58 4003
rect 52 3998 53 4002
rect 57 3998 58 4002
rect 111 4000 112 4004
rect 116 4000 119 4004
rect 123 4000 125 4004
rect 129 4000 131 4004
rect 107 3998 135 4000
rect 4 3994 14 3998
rect 18 3994 20 3998
rect 24 3994 26 3998
rect 30 3994 32 3998
rect 36 3994 38 3998
rect 42 3994 43 3998
rect 47 3994 48 3998
rect 111 3994 112 3998
rect 116 3994 119 3998
rect 123 3994 125 3998
rect 129 3994 131 3998
rect 0 3993 100 3994
rect 0 3992 64 3993
rect 4 3988 14 3992
rect 18 3988 20 3992
rect 24 3988 26 3992
rect 30 3988 32 3992
rect 36 3988 38 3992
rect 42 3988 43 3992
rect 47 3989 64 3992
rect 68 3989 70 3993
rect 74 3989 76 3993
rect 80 3989 82 3993
rect 86 3989 89 3993
rect 93 3989 95 3993
rect 99 3989 100 3993
rect 47 3988 100 3989
rect 0 3987 100 3988
rect 0 3986 64 3987
rect 4 3982 14 3986
rect 18 3982 20 3986
rect 24 3982 26 3986
rect 30 3982 32 3986
rect 36 3982 38 3986
rect 42 3982 43 3986
rect 47 3983 64 3986
rect 68 3983 70 3987
rect 74 3983 76 3987
rect 80 3983 82 3987
rect 86 3983 89 3987
rect 93 3983 95 3987
rect 99 3983 100 3987
rect 47 3982 100 3983
rect 0 3981 100 3982
rect 0 3980 64 3981
rect 4 3976 14 3980
rect 18 3976 20 3980
rect 24 3976 26 3980
rect 30 3976 32 3980
rect 36 3976 38 3980
rect 42 3976 43 3980
rect 47 3977 64 3980
rect 68 3977 70 3981
rect 74 3977 76 3981
rect 80 3977 82 3981
rect 86 3977 89 3981
rect 93 3977 95 3981
rect 99 3977 100 3981
rect 47 3976 100 3977
rect 0 3975 100 3976
rect 0 3974 64 3975
rect 4 3970 14 3974
rect 18 3970 20 3974
rect 24 3970 26 3974
rect 30 3970 32 3974
rect 36 3970 38 3974
rect 42 3970 43 3974
rect 47 3971 64 3974
rect 68 3971 70 3975
rect 74 3971 76 3975
rect 80 3971 82 3975
rect 86 3971 89 3975
rect 93 3971 95 3975
rect 99 3971 100 3975
rect 47 3970 100 3971
rect 0 3969 100 3970
rect 0 3968 64 3969
rect 4 3964 20 3968
rect 24 3964 26 3968
rect 30 3964 32 3968
rect 36 3964 38 3968
rect 42 3964 43 3968
rect 47 3965 64 3968
rect 68 3965 70 3969
rect 74 3965 76 3969
rect 80 3965 82 3969
rect 86 3965 89 3969
rect 93 3965 95 3969
rect 99 3965 100 3969
rect 47 3964 100 3965
rect 107 3992 135 3994
rect 111 3988 112 3992
rect 116 3988 119 3992
rect 123 3988 125 3992
rect 129 3988 131 3992
rect 107 3986 135 3988
rect 111 3982 112 3986
rect 116 3982 119 3986
rect 123 3982 125 3986
rect 129 3982 131 3986
rect 107 3980 135 3982
rect 111 3976 112 3980
rect 116 3976 119 3980
rect 123 3976 125 3980
rect 129 3976 131 3980
rect 107 3974 135 3976
rect 111 3970 112 3974
rect 116 3970 119 3974
rect 123 3970 125 3974
rect 129 3970 131 3974
rect 144 3998 148 4000
rect 144 3992 148 3994
rect 144 3986 148 3988
rect 144 3980 148 3982
rect 144 3974 148 3976
rect 107 3968 129 3970
rect 111 3964 112 3968
rect 116 3964 119 3968
rect 123 3964 125 3968
rect 144 3968 148 3970
rect 144 3962 148 3964
rect 4 3956 8 3960
rect 12 3956 63 3960
rect 72 3956 74 3960
rect 78 3956 80 3960
rect 84 3956 86 3960
rect 90 3956 92 3960
rect 101 3956 137 3960
rect 141 3958 144 3960
rect 141 3956 148 3958
rect 0 3954 144 3956
rect 4 3950 8 3954
rect 12 3950 63 3954
rect 72 3950 74 3954
rect 78 3950 80 3954
rect 84 3950 86 3954
rect 90 3950 92 3954
rect 101 3950 137 3954
rect 141 3952 144 3954
rect 141 3950 148 3952
rect 0 3948 144 3950
rect 4 3944 8 3948
rect 12 3944 63 3948
rect 72 3944 74 3948
rect 78 3944 80 3948
rect 84 3944 86 3948
rect 90 3944 92 3948
rect 101 3944 137 3948
rect 141 3946 144 3948
rect 141 3944 148 3946
rect 0 3942 144 3944
rect 4 3938 8 3942
rect 12 3938 63 3942
rect 72 3938 74 3942
rect 78 3938 80 3942
rect 84 3938 86 3942
rect 90 3938 92 3942
rect 101 3938 137 3942
rect 141 3940 144 3942
rect 141 3938 148 3940
rect 0 3936 144 3938
rect 4 3932 8 3936
rect 12 3932 63 3936
rect 72 3932 74 3936
rect 78 3932 80 3936
rect 84 3932 86 3936
rect 90 3932 92 3936
rect 101 3932 137 3936
rect 141 3934 144 3936
rect 141 3932 148 3934
rect 0 3930 144 3932
rect 4 3926 8 3930
rect 12 3926 63 3930
rect 72 3926 74 3930
rect 78 3926 80 3930
rect 84 3926 86 3930
rect 90 3926 92 3930
rect 101 3926 137 3930
rect 141 3928 144 3930
rect 141 3926 148 3928
rect 0 3924 144 3926
rect 4 3920 8 3924
rect 12 3920 63 3924
rect 72 3920 74 3924
rect 78 3920 80 3924
rect 84 3920 86 3924
rect 90 3920 92 3924
rect 101 3920 137 3924
rect 141 3922 144 3924
rect 141 3920 148 3922
rect 144 3914 148 3916
rect 144 3908 148 3910
rect 144 3902 148 3904
rect 144 3896 148 3898
rect 144 3890 148 3892
rect 144 3884 148 3886
rect 144 3878 148 3880
rect 144 3872 148 3874
rect 144 3866 148 3868
rect 144 3860 148 3862
rect 144 3854 148 3856
rect 144 3848 148 3850
rect 144 3842 148 3844
rect 144 3836 148 3838
rect 144 3830 148 3832
rect 144 3824 148 3826
rect 144 3818 148 3820
rect 144 3812 148 3814
rect 144 3806 148 3808
rect 144 3800 148 3802
rect 144 3794 148 3796
rect 148 3790 150 3794
rect 154 3790 156 3794
rect 160 3790 162 3794
rect 166 3790 168 3794
rect 172 3790 174 3794
rect 178 3790 180 3794
rect 184 3790 186 3794
rect 190 3790 192 3794
rect 196 3790 198 3794
rect 202 3790 204 3794
rect 208 3790 210 3794
rect 214 3790 216 3794
rect 220 3790 222 3794
rect 226 3790 228 3794
rect 232 3790 234 3794
rect 238 3790 240 3794
rect 244 3790 246 3794
rect 250 3790 252 3794
rect 256 3790 258 3794
rect 262 3790 264 3794
rect 268 3790 270 3794
rect 274 3790 276 3794
rect 280 3790 282 3794
rect 286 3790 288 3794
rect 292 3790 294 3794
rect 298 3790 300 3794
rect 304 3790 306 3794
rect 310 3790 312 3794
rect 316 3790 318 3794
rect 322 3790 324 3794
rect 328 3790 330 3794
rect 334 3790 336 3794
rect 340 3790 342 3794
rect 346 3790 348 3794
rect 352 3790 354 3794
rect 358 3790 360 3794
rect 364 3790 366 3794
rect 370 3790 372 3794
rect 376 3790 378 3794
rect 382 3790 384 3794
rect 388 3790 390 3794
rect 394 3790 396 3794
rect 400 3790 402 3794
rect 406 3790 408 3794
rect 412 3790 414 3794
rect 418 3790 420 3794
rect 424 3790 426 3794
rect 430 3790 432 3794
rect 436 3790 438 3794
rect 442 3790 444 3794
rect 448 3790 450 3794
rect 454 3790 456 3794
rect 460 3790 462 3794
rect 466 3790 468 3794
rect 472 3790 474 3794
rect 478 3790 480 3794
rect 484 3790 486 3794
rect 490 3790 492 3794
rect 496 3790 498 3794
rect 502 3790 504 3794
rect 508 3790 510 3794
rect 144 3788 148 3790
rect 144 3782 148 3784
rect 144 3776 148 3778
rect 144 3770 148 3772
rect 144 3764 148 3766
rect 144 3758 148 3760
rect 144 3752 148 3754
rect 144 3746 148 3748
rect 144 3740 148 3742
rect 144 3734 148 3736
rect 144 3728 148 3730
rect 144 3722 148 3724
rect 144 3716 148 3718
rect 144 3710 148 3712
rect 144 3704 148 3706
rect 144 3698 148 3700
rect 144 3692 148 3694
rect 144 3686 148 3688
rect 144 3680 148 3682
rect 144 3674 148 3676
rect 144 3668 148 3670
rect 4 3660 8 3664
rect 12 3660 63 3664
rect 72 3660 74 3664
rect 78 3660 80 3664
rect 84 3660 86 3664
rect 90 3660 92 3664
rect 101 3660 137 3664
rect 141 3662 148 3664
rect 141 3660 144 3662
rect 0 3658 144 3660
rect 4 3654 8 3658
rect 12 3654 63 3658
rect 72 3654 74 3658
rect 78 3654 80 3658
rect 84 3654 86 3658
rect 90 3654 92 3658
rect 101 3654 137 3658
rect 141 3656 148 3658
rect 141 3654 144 3656
rect 0 3652 144 3654
rect 4 3648 8 3652
rect 12 3648 63 3652
rect 72 3648 74 3652
rect 78 3648 80 3652
rect 84 3648 86 3652
rect 90 3648 92 3652
rect 101 3648 137 3652
rect 141 3650 148 3652
rect 141 3648 144 3650
rect 0 3646 144 3648
rect 4 3642 8 3646
rect 12 3642 63 3646
rect 72 3642 74 3646
rect 78 3642 80 3646
rect 84 3642 86 3646
rect 90 3642 92 3646
rect 101 3642 137 3646
rect 141 3644 148 3646
rect 141 3642 144 3644
rect 0 3640 144 3642
rect 4 3636 8 3640
rect 12 3636 63 3640
rect 72 3636 74 3640
rect 78 3636 80 3640
rect 84 3636 86 3640
rect 90 3636 92 3640
rect 101 3636 137 3640
rect 141 3638 148 3640
rect 141 3636 144 3638
rect 0 3634 144 3636
rect 4 3630 8 3634
rect 12 3630 63 3634
rect 72 3630 74 3634
rect 78 3630 80 3634
rect 84 3630 86 3634
rect 90 3630 92 3634
rect 101 3630 137 3634
rect 141 3632 148 3634
rect 141 3630 144 3632
rect 0 3628 144 3630
rect 4 3624 8 3628
rect 12 3624 63 3628
rect 72 3624 74 3628
rect 78 3624 80 3628
rect 84 3624 86 3628
rect 90 3624 92 3628
rect 101 3624 137 3628
rect 141 3626 148 3628
rect 141 3624 144 3626
rect 144 3620 148 3622
rect 4 3616 20 3620
rect 24 3616 26 3620
rect 30 3616 32 3620
rect 36 3616 38 3620
rect 42 3616 44 3620
rect 48 3619 100 3620
rect 48 3616 64 3619
rect 0 3615 64 3616
rect 68 3615 70 3619
rect 74 3615 76 3619
rect 80 3615 82 3619
rect 86 3615 89 3619
rect 93 3615 95 3619
rect 99 3615 100 3619
rect 0 3614 100 3615
rect 4 3610 14 3614
rect 18 3610 20 3614
rect 24 3610 26 3614
rect 30 3610 32 3614
rect 36 3610 38 3614
rect 42 3610 44 3614
rect 48 3613 100 3614
rect 48 3610 64 3613
rect 0 3609 64 3610
rect 68 3609 70 3613
rect 74 3609 76 3613
rect 80 3609 82 3613
rect 86 3609 89 3613
rect 93 3609 95 3613
rect 99 3609 100 3613
rect 0 3608 100 3609
rect 4 3604 14 3608
rect 18 3604 20 3608
rect 24 3604 26 3608
rect 30 3604 32 3608
rect 36 3604 38 3608
rect 42 3604 44 3608
rect 48 3607 100 3608
rect 48 3604 64 3607
rect 0 3603 64 3604
rect 68 3603 70 3607
rect 74 3603 76 3607
rect 80 3603 82 3607
rect 86 3603 89 3607
rect 93 3603 95 3607
rect 99 3603 100 3607
rect 0 3602 100 3603
rect 4 3598 14 3602
rect 18 3598 20 3602
rect 24 3598 26 3602
rect 30 3598 32 3602
rect 36 3598 38 3602
rect 42 3598 44 3602
rect 48 3601 100 3602
rect 48 3598 64 3601
rect 0 3597 64 3598
rect 68 3597 70 3601
rect 74 3597 76 3601
rect 80 3597 82 3601
rect 86 3597 89 3601
rect 93 3597 95 3601
rect 99 3597 100 3601
rect 0 3596 100 3597
rect 4 3592 14 3596
rect 18 3592 20 3596
rect 24 3592 26 3596
rect 30 3592 32 3596
rect 36 3592 38 3596
rect 42 3592 44 3596
rect 48 3595 100 3596
rect 48 3592 64 3595
rect 0 3591 64 3592
rect 68 3591 70 3595
rect 74 3591 76 3595
rect 80 3591 82 3595
rect 86 3591 89 3595
rect 93 3591 95 3595
rect 99 3591 100 3595
rect 0 3590 100 3591
rect 111 3616 112 3620
rect 116 3616 119 3620
rect 123 3616 125 3620
rect 107 3614 129 3616
rect 144 3614 148 3616
rect 111 3610 112 3614
rect 116 3610 119 3614
rect 123 3610 125 3614
rect 129 3610 131 3614
rect 107 3608 135 3610
rect 111 3604 112 3608
rect 116 3604 119 3608
rect 123 3604 125 3608
rect 129 3604 131 3608
rect 107 3602 135 3604
rect 111 3598 112 3602
rect 116 3598 119 3602
rect 123 3598 125 3602
rect 129 3598 131 3602
rect 107 3596 135 3598
rect 111 3592 112 3596
rect 116 3592 119 3596
rect 123 3592 125 3596
rect 129 3592 131 3596
rect 107 3590 135 3592
rect 4 3586 14 3590
rect 18 3586 20 3590
rect 24 3586 26 3590
rect 30 3586 32 3590
rect 36 3586 38 3590
rect 42 3586 44 3590
rect 111 3586 112 3590
rect 116 3586 119 3590
rect 123 3586 125 3590
rect 129 3586 131 3590
rect 0 3584 48 3586
rect 4 3580 14 3584
rect 18 3580 20 3584
rect 24 3580 26 3584
rect 30 3580 32 3584
rect 36 3580 38 3584
rect 42 3580 44 3584
rect 52 3582 53 3586
rect 57 3582 58 3586
rect 52 3581 58 3582
rect 52 3577 53 3581
rect 57 3577 58 3581
rect 107 3584 135 3586
rect 111 3580 112 3584
rect 116 3580 119 3584
rect 123 3580 125 3584
rect 129 3580 131 3584
rect 144 3608 148 3610
rect 144 3602 148 3604
rect 144 3596 148 3598
rect 144 3590 148 3592
rect 144 3584 148 3586
rect 52 3576 58 3577
rect 4 3572 53 3576
rect 57 3572 58 3576
rect 4 3571 58 3572
rect 4 3567 53 3571
rect 57 3567 58 3571
rect 144 3578 148 3580
rect 144 3572 148 3574
rect 4 3539 53 3543
rect 57 3539 58 3543
rect 4 3538 58 3539
rect 4 3534 53 3538
rect 57 3534 58 3538
rect 52 3533 58 3534
rect 4 3526 14 3530
rect 18 3526 20 3530
rect 24 3526 26 3530
rect 30 3526 32 3530
rect 36 3526 38 3530
rect 42 3526 44 3530
rect 0 3524 48 3526
rect 52 3529 53 3533
rect 57 3529 58 3533
rect 144 3536 148 3538
rect 144 3530 148 3532
rect 52 3528 58 3529
rect 52 3524 53 3528
rect 57 3524 58 3528
rect 111 3526 112 3530
rect 116 3526 119 3530
rect 123 3526 125 3530
rect 129 3526 131 3530
rect 107 3524 135 3526
rect 4 3520 14 3524
rect 18 3520 20 3524
rect 24 3520 26 3524
rect 30 3520 32 3524
rect 36 3520 38 3524
rect 42 3520 44 3524
rect 111 3520 112 3524
rect 116 3520 119 3524
rect 123 3520 125 3524
rect 129 3520 131 3524
rect 0 3519 100 3520
rect 0 3518 64 3519
rect 4 3514 14 3518
rect 18 3514 20 3518
rect 24 3514 26 3518
rect 30 3514 32 3518
rect 36 3514 38 3518
rect 42 3514 44 3518
rect 48 3515 64 3518
rect 68 3515 70 3519
rect 74 3515 76 3519
rect 80 3515 82 3519
rect 86 3515 89 3519
rect 93 3515 95 3519
rect 99 3515 100 3519
rect 48 3514 100 3515
rect 0 3513 100 3514
rect 0 3512 64 3513
rect 4 3508 14 3512
rect 18 3508 20 3512
rect 24 3508 26 3512
rect 30 3508 32 3512
rect 36 3508 38 3512
rect 42 3508 44 3512
rect 48 3509 64 3512
rect 68 3509 70 3513
rect 74 3509 76 3513
rect 80 3509 82 3513
rect 86 3509 89 3513
rect 93 3509 95 3513
rect 99 3509 100 3513
rect 48 3508 100 3509
rect 0 3507 100 3508
rect 0 3506 64 3507
rect 4 3502 14 3506
rect 18 3502 20 3506
rect 24 3502 26 3506
rect 30 3502 32 3506
rect 36 3502 38 3506
rect 42 3502 44 3506
rect 48 3503 64 3506
rect 68 3503 70 3507
rect 74 3503 76 3507
rect 80 3503 82 3507
rect 86 3503 89 3507
rect 93 3503 95 3507
rect 99 3503 100 3507
rect 48 3502 100 3503
rect 0 3501 100 3502
rect 0 3500 64 3501
rect 4 3496 14 3500
rect 18 3496 20 3500
rect 24 3496 26 3500
rect 30 3496 32 3500
rect 36 3496 38 3500
rect 42 3496 44 3500
rect 48 3497 64 3500
rect 68 3497 70 3501
rect 74 3497 76 3501
rect 80 3497 82 3501
rect 86 3497 89 3501
rect 93 3497 95 3501
rect 99 3497 100 3501
rect 48 3496 100 3497
rect 0 3495 100 3496
rect 0 3494 64 3495
rect 4 3490 20 3494
rect 24 3490 26 3494
rect 30 3490 32 3494
rect 36 3490 38 3494
rect 42 3490 44 3494
rect 48 3491 64 3494
rect 68 3491 70 3495
rect 74 3491 76 3495
rect 80 3491 82 3495
rect 86 3491 89 3495
rect 93 3491 95 3495
rect 99 3491 100 3495
rect 48 3490 100 3491
rect 107 3518 135 3520
rect 111 3514 112 3518
rect 116 3514 119 3518
rect 123 3514 125 3518
rect 129 3514 131 3518
rect 107 3512 135 3514
rect 111 3508 112 3512
rect 116 3508 119 3512
rect 123 3508 125 3512
rect 129 3508 131 3512
rect 107 3506 135 3508
rect 111 3502 112 3506
rect 116 3502 119 3506
rect 123 3502 125 3506
rect 129 3502 131 3506
rect 107 3500 135 3502
rect 111 3496 112 3500
rect 116 3496 119 3500
rect 123 3496 125 3500
rect 129 3496 131 3500
rect 144 3524 148 3526
rect 144 3518 148 3520
rect 144 3512 148 3514
rect 144 3506 148 3508
rect 144 3500 148 3502
rect 107 3494 129 3496
rect 111 3490 112 3494
rect 116 3490 119 3494
rect 123 3490 125 3494
rect 144 3494 148 3496
rect 144 3488 148 3490
rect 4 3482 8 3486
rect 12 3482 63 3486
rect 72 3482 74 3486
rect 78 3482 80 3486
rect 84 3482 86 3486
rect 90 3482 92 3486
rect 101 3482 137 3486
rect 141 3484 144 3486
rect 141 3482 148 3484
rect 0 3480 144 3482
rect 4 3476 8 3480
rect 12 3476 63 3480
rect 72 3476 74 3480
rect 78 3476 80 3480
rect 84 3476 86 3480
rect 90 3476 92 3480
rect 101 3476 137 3480
rect 141 3478 144 3480
rect 141 3476 148 3478
rect 0 3474 144 3476
rect 4 3470 8 3474
rect 12 3470 63 3474
rect 72 3470 74 3474
rect 78 3470 80 3474
rect 84 3470 86 3474
rect 90 3470 92 3474
rect 101 3470 137 3474
rect 141 3472 144 3474
rect 141 3470 148 3472
rect 0 3468 144 3470
rect 4 3464 8 3468
rect 12 3464 63 3468
rect 72 3464 74 3468
rect 78 3464 80 3468
rect 84 3464 86 3468
rect 90 3464 92 3468
rect 101 3464 137 3468
rect 141 3466 144 3468
rect 141 3464 148 3466
rect 0 3462 144 3464
rect 4 3458 8 3462
rect 12 3458 63 3462
rect 72 3458 74 3462
rect 78 3458 80 3462
rect 84 3458 86 3462
rect 90 3458 92 3462
rect 101 3458 137 3462
rect 141 3460 144 3462
rect 141 3458 148 3460
rect 0 3456 144 3458
rect 4 3452 8 3456
rect 12 3452 63 3456
rect 72 3452 74 3456
rect 78 3452 80 3456
rect 84 3452 86 3456
rect 90 3452 92 3456
rect 101 3452 137 3456
rect 141 3454 144 3456
rect 141 3452 148 3454
rect 0 3450 144 3452
rect 4 3446 8 3450
rect 12 3446 63 3450
rect 72 3446 74 3450
rect 78 3446 80 3450
rect 84 3446 86 3450
rect 90 3446 92 3450
rect 101 3446 137 3450
rect 141 3448 144 3450
rect 141 3446 148 3448
rect 144 3440 148 3442
rect 144 3434 148 3436
rect 144 3428 148 3430
rect 144 3422 148 3424
rect 144 3416 148 3418
rect 144 3410 148 3412
rect 144 3404 148 3406
rect 144 3398 148 3400
rect 144 3392 148 3394
rect 144 3386 148 3388
rect 144 3380 148 3382
rect 144 3374 148 3376
rect 144 3368 148 3370
rect 144 3362 148 3364
rect 144 3356 148 3358
rect 144 3350 148 3352
rect 144 3344 148 3346
rect 144 3338 148 3340
rect 144 3332 148 3334
rect 144 3326 148 3328
rect 144 3320 148 3322
rect 148 3316 150 3320
rect 154 3316 156 3320
rect 160 3316 162 3320
rect 166 3316 168 3320
rect 172 3316 174 3320
rect 178 3316 180 3320
rect 184 3316 186 3320
rect 190 3316 192 3320
rect 196 3316 198 3320
rect 202 3316 204 3320
rect 208 3316 210 3320
rect 214 3316 216 3320
rect 220 3316 222 3320
rect 226 3316 228 3320
rect 232 3316 234 3320
rect 238 3316 240 3320
rect 244 3316 246 3320
rect 250 3316 252 3320
rect 256 3316 258 3320
rect 262 3316 264 3320
rect 268 3316 270 3320
rect 274 3316 276 3320
rect 280 3316 282 3320
rect 286 3316 288 3320
rect 292 3316 294 3320
rect 298 3316 300 3320
rect 304 3316 306 3320
rect 310 3316 312 3320
rect 316 3316 318 3320
rect 322 3316 324 3320
rect 328 3316 330 3320
rect 334 3316 336 3320
rect 340 3316 342 3320
rect 346 3316 348 3320
rect 352 3316 354 3320
rect 358 3316 360 3320
rect 364 3316 366 3320
rect 370 3316 372 3320
rect 376 3316 378 3320
rect 382 3316 384 3320
rect 388 3316 390 3320
rect 394 3316 396 3320
rect 400 3316 402 3320
rect 406 3316 408 3320
rect 412 3316 414 3320
rect 418 3316 420 3320
rect 424 3316 426 3320
rect 430 3316 432 3320
rect 436 3316 438 3320
rect 442 3316 444 3320
rect 448 3316 450 3320
rect 454 3316 456 3320
rect 460 3316 462 3320
rect 466 3316 468 3320
rect 472 3316 474 3320
rect 478 3316 480 3320
rect 484 3316 486 3320
rect 490 3316 492 3320
rect 496 3316 498 3320
rect 502 3316 504 3320
rect 508 3316 510 3320
rect 144 3314 148 3316
rect 144 3308 148 3310
rect 144 3302 148 3304
rect 144 3296 148 3298
rect 144 3290 148 3292
rect 144 3284 148 3286
rect 144 3278 148 3280
rect 144 3272 148 3274
rect 144 3266 148 3268
rect 144 3260 148 3262
rect 144 3254 148 3256
rect 144 3248 148 3250
rect 144 3242 148 3244
rect 144 3236 148 3238
rect 144 3230 148 3232
rect 144 3224 148 3226
rect 144 3218 148 3220
rect 144 3212 148 3214
rect 144 3206 148 3208
rect 144 3200 148 3202
rect 144 3194 148 3196
rect 4 3186 8 3190
rect 12 3186 63 3190
rect 72 3186 74 3190
rect 78 3186 80 3190
rect 84 3186 86 3190
rect 90 3186 92 3190
rect 101 3186 137 3190
rect 141 3188 148 3190
rect 141 3186 144 3188
rect 0 3184 144 3186
rect 4 3180 8 3184
rect 12 3180 63 3184
rect 72 3180 74 3184
rect 78 3180 80 3184
rect 84 3180 86 3184
rect 90 3180 92 3184
rect 101 3180 137 3184
rect 141 3182 148 3184
rect 141 3180 144 3182
rect 0 3178 144 3180
rect 4 3174 8 3178
rect 12 3174 63 3178
rect 72 3174 74 3178
rect 78 3174 80 3178
rect 84 3174 86 3178
rect 90 3174 92 3178
rect 101 3174 137 3178
rect 141 3176 148 3178
rect 141 3174 144 3176
rect 0 3172 144 3174
rect 4 3168 8 3172
rect 12 3168 63 3172
rect 72 3168 74 3172
rect 78 3168 80 3172
rect 84 3168 86 3172
rect 90 3168 92 3172
rect 101 3168 137 3172
rect 141 3170 148 3172
rect 141 3168 144 3170
rect 0 3166 144 3168
rect 4 3162 8 3166
rect 12 3162 63 3166
rect 72 3162 74 3166
rect 78 3162 80 3166
rect 84 3162 86 3166
rect 90 3162 92 3166
rect 101 3162 137 3166
rect 141 3164 148 3166
rect 141 3162 144 3164
rect 0 3160 144 3162
rect 4 3156 8 3160
rect 12 3156 63 3160
rect 72 3156 74 3160
rect 78 3156 80 3160
rect 84 3156 86 3160
rect 90 3156 92 3160
rect 101 3156 137 3160
rect 141 3158 148 3160
rect 141 3156 144 3158
rect 0 3154 144 3156
rect 4 3150 8 3154
rect 12 3150 63 3154
rect 72 3150 74 3154
rect 78 3150 80 3154
rect 84 3150 86 3154
rect 90 3150 92 3154
rect 101 3150 137 3154
rect 141 3152 148 3154
rect 141 3150 144 3152
rect 144 3146 148 3148
rect 4 3142 20 3146
rect 24 3142 26 3146
rect 30 3142 32 3146
rect 36 3142 38 3146
rect 42 3142 44 3146
rect 48 3145 100 3146
rect 48 3142 64 3145
rect 0 3141 64 3142
rect 68 3141 70 3145
rect 74 3141 76 3145
rect 80 3141 82 3145
rect 86 3141 89 3145
rect 93 3141 95 3145
rect 99 3141 100 3145
rect 0 3140 100 3141
rect 4 3136 14 3140
rect 18 3136 20 3140
rect 24 3136 26 3140
rect 30 3136 32 3140
rect 36 3136 38 3140
rect 42 3136 44 3140
rect 48 3139 100 3140
rect 48 3136 64 3139
rect 0 3135 64 3136
rect 68 3135 70 3139
rect 74 3135 76 3139
rect 80 3135 82 3139
rect 86 3135 89 3139
rect 93 3135 95 3139
rect 99 3135 100 3139
rect 0 3134 100 3135
rect 4 3130 14 3134
rect 18 3130 20 3134
rect 24 3130 26 3134
rect 30 3130 32 3134
rect 36 3130 38 3134
rect 42 3130 44 3134
rect 48 3133 100 3134
rect 48 3130 64 3133
rect 0 3129 64 3130
rect 68 3129 70 3133
rect 74 3129 76 3133
rect 80 3129 82 3133
rect 86 3129 89 3133
rect 93 3129 95 3133
rect 99 3129 100 3133
rect 0 3128 100 3129
rect 4 3124 14 3128
rect 18 3124 20 3128
rect 24 3124 26 3128
rect 30 3124 32 3128
rect 36 3124 38 3128
rect 42 3124 44 3128
rect 48 3127 100 3128
rect 48 3124 64 3127
rect 0 3123 64 3124
rect 68 3123 70 3127
rect 74 3123 76 3127
rect 80 3123 82 3127
rect 86 3123 89 3127
rect 93 3123 95 3127
rect 99 3123 100 3127
rect 0 3122 100 3123
rect 4 3118 14 3122
rect 18 3118 20 3122
rect 24 3118 26 3122
rect 30 3118 32 3122
rect 36 3118 38 3122
rect 42 3118 44 3122
rect 48 3121 100 3122
rect 48 3118 64 3121
rect 0 3117 64 3118
rect 68 3117 70 3121
rect 74 3117 76 3121
rect 80 3117 82 3121
rect 86 3117 89 3121
rect 93 3117 95 3121
rect 99 3117 100 3121
rect 0 3116 100 3117
rect 111 3142 112 3146
rect 116 3142 119 3146
rect 123 3142 125 3146
rect 107 3140 129 3142
rect 144 3140 148 3142
rect 111 3136 112 3140
rect 116 3136 119 3140
rect 123 3136 125 3140
rect 129 3136 131 3140
rect 107 3134 135 3136
rect 111 3130 112 3134
rect 116 3130 119 3134
rect 123 3130 125 3134
rect 129 3130 131 3134
rect 107 3128 135 3130
rect 111 3124 112 3128
rect 116 3124 119 3128
rect 123 3124 125 3128
rect 129 3124 131 3128
rect 107 3122 135 3124
rect 111 3118 112 3122
rect 116 3118 119 3122
rect 123 3118 125 3122
rect 129 3118 131 3122
rect 107 3116 135 3118
rect 4 3112 14 3116
rect 18 3112 20 3116
rect 24 3112 26 3116
rect 30 3112 32 3116
rect 36 3112 38 3116
rect 42 3112 44 3116
rect 111 3112 112 3116
rect 116 3112 119 3116
rect 123 3112 125 3116
rect 129 3112 131 3116
rect 0 3110 48 3112
rect 4 3106 14 3110
rect 18 3106 20 3110
rect 24 3106 26 3110
rect 30 3106 32 3110
rect 36 3106 38 3110
rect 42 3106 44 3110
rect 52 3108 53 3112
rect 57 3108 58 3112
rect 52 3107 58 3108
rect 52 3103 53 3107
rect 57 3103 58 3107
rect 107 3110 135 3112
rect 111 3106 112 3110
rect 116 3106 119 3110
rect 123 3106 125 3110
rect 129 3106 131 3110
rect 144 3134 148 3136
rect 144 3128 148 3130
rect 144 3122 148 3124
rect 144 3116 148 3118
rect 144 3110 148 3112
rect 52 3102 58 3103
rect 4 3098 53 3102
rect 57 3098 58 3102
rect 4 3097 58 3098
rect 4 3093 53 3097
rect 57 3093 58 3097
rect 144 3104 148 3106
rect 144 3098 148 3100
rect 4 3065 53 3069
rect 57 3065 58 3069
rect 4 3064 58 3065
rect 4 3060 53 3064
rect 57 3060 58 3064
rect 52 3059 58 3060
rect 4 3052 14 3056
rect 18 3052 20 3056
rect 24 3052 26 3056
rect 30 3052 32 3056
rect 36 3052 38 3056
rect 42 3052 44 3056
rect 0 3050 48 3052
rect 52 3055 53 3059
rect 57 3055 58 3059
rect 144 3062 148 3064
rect 144 3056 148 3058
rect 52 3054 58 3055
rect 52 3050 53 3054
rect 57 3050 58 3054
rect 111 3052 112 3056
rect 116 3052 119 3056
rect 123 3052 125 3056
rect 129 3052 131 3056
rect 107 3050 135 3052
rect 4 3046 14 3050
rect 18 3046 20 3050
rect 24 3046 26 3050
rect 30 3046 32 3050
rect 36 3046 38 3050
rect 42 3046 44 3050
rect 111 3046 112 3050
rect 116 3046 119 3050
rect 123 3046 125 3050
rect 129 3046 131 3050
rect 0 3045 100 3046
rect 0 3044 64 3045
rect 4 3040 14 3044
rect 18 3040 20 3044
rect 24 3040 26 3044
rect 30 3040 32 3044
rect 36 3040 38 3044
rect 42 3040 44 3044
rect 48 3041 64 3044
rect 68 3041 70 3045
rect 74 3041 76 3045
rect 80 3041 82 3045
rect 86 3041 89 3045
rect 93 3041 95 3045
rect 99 3041 100 3045
rect 48 3040 100 3041
rect 0 3039 100 3040
rect 0 3038 64 3039
rect 4 3034 14 3038
rect 18 3034 20 3038
rect 24 3034 26 3038
rect 30 3034 32 3038
rect 36 3034 38 3038
rect 42 3034 44 3038
rect 48 3035 64 3038
rect 68 3035 70 3039
rect 74 3035 76 3039
rect 80 3035 82 3039
rect 86 3035 89 3039
rect 93 3035 95 3039
rect 99 3035 100 3039
rect 48 3034 100 3035
rect 0 3033 100 3034
rect 0 3032 64 3033
rect 4 3028 14 3032
rect 18 3028 20 3032
rect 24 3028 26 3032
rect 30 3028 32 3032
rect 36 3028 38 3032
rect 42 3028 44 3032
rect 48 3029 64 3032
rect 68 3029 70 3033
rect 74 3029 76 3033
rect 80 3029 82 3033
rect 86 3029 89 3033
rect 93 3029 95 3033
rect 99 3029 100 3033
rect 48 3028 100 3029
rect 0 3027 100 3028
rect 0 3026 64 3027
rect 4 3022 14 3026
rect 18 3022 20 3026
rect 24 3022 26 3026
rect 30 3022 32 3026
rect 36 3022 38 3026
rect 42 3022 44 3026
rect 48 3023 64 3026
rect 68 3023 70 3027
rect 74 3023 76 3027
rect 80 3023 82 3027
rect 86 3023 89 3027
rect 93 3023 95 3027
rect 99 3023 100 3027
rect 48 3022 100 3023
rect 0 3021 100 3022
rect 0 3020 64 3021
rect 4 3016 20 3020
rect 24 3016 26 3020
rect 30 3016 32 3020
rect 36 3016 38 3020
rect 42 3016 44 3020
rect 48 3017 64 3020
rect 68 3017 70 3021
rect 74 3017 76 3021
rect 80 3017 82 3021
rect 86 3017 89 3021
rect 93 3017 95 3021
rect 99 3017 100 3021
rect 48 3016 100 3017
rect 107 3044 135 3046
rect 111 3040 112 3044
rect 116 3040 119 3044
rect 123 3040 125 3044
rect 129 3040 131 3044
rect 107 3038 135 3040
rect 111 3034 112 3038
rect 116 3034 119 3038
rect 123 3034 125 3038
rect 129 3034 131 3038
rect 107 3032 135 3034
rect 111 3028 112 3032
rect 116 3028 119 3032
rect 123 3028 125 3032
rect 129 3028 131 3032
rect 107 3026 135 3028
rect 111 3022 112 3026
rect 116 3022 119 3026
rect 123 3022 125 3026
rect 129 3022 131 3026
rect 144 3050 148 3052
rect 144 3044 148 3046
rect 144 3038 148 3040
rect 144 3032 148 3034
rect 144 3026 148 3028
rect 107 3020 129 3022
rect 111 3016 112 3020
rect 116 3016 119 3020
rect 123 3016 125 3020
rect 144 3020 148 3022
rect 144 3014 148 3016
rect 4 3008 8 3012
rect 12 3008 63 3012
rect 72 3008 74 3012
rect 78 3008 80 3012
rect 84 3008 86 3012
rect 90 3008 92 3012
rect 101 3008 137 3012
rect 141 3010 144 3012
rect 141 3008 148 3010
rect 0 3006 144 3008
rect 4 3002 8 3006
rect 12 3002 63 3006
rect 72 3002 74 3006
rect 78 3002 80 3006
rect 84 3002 86 3006
rect 90 3002 92 3006
rect 101 3002 137 3006
rect 141 3004 144 3006
rect 141 3002 148 3004
rect 0 3000 144 3002
rect 4 2996 8 3000
rect 12 2996 63 3000
rect 72 2996 74 3000
rect 78 2996 80 3000
rect 84 2996 86 3000
rect 90 2996 92 3000
rect 101 2996 137 3000
rect 141 2998 144 3000
rect 141 2996 148 2998
rect 0 2994 144 2996
rect 4 2990 8 2994
rect 12 2990 63 2994
rect 72 2990 74 2994
rect 78 2990 80 2994
rect 84 2990 86 2994
rect 90 2990 92 2994
rect 101 2990 137 2994
rect 141 2992 144 2994
rect 141 2990 148 2992
rect 0 2988 144 2990
rect 4 2984 8 2988
rect 12 2984 63 2988
rect 72 2984 74 2988
rect 78 2984 80 2988
rect 84 2984 86 2988
rect 90 2984 92 2988
rect 101 2984 137 2988
rect 141 2986 144 2988
rect 141 2984 148 2986
rect 0 2982 144 2984
rect 4 2978 8 2982
rect 12 2978 63 2982
rect 72 2978 74 2982
rect 78 2978 80 2982
rect 84 2978 86 2982
rect 90 2978 92 2982
rect 101 2978 137 2982
rect 141 2980 144 2982
rect 141 2978 148 2980
rect 0 2976 144 2978
rect 4 2972 8 2976
rect 12 2972 63 2976
rect 72 2972 74 2976
rect 78 2972 80 2976
rect 84 2972 86 2976
rect 90 2972 92 2976
rect 101 2972 137 2976
rect 141 2974 144 2976
rect 141 2972 148 2974
rect 144 2966 148 2968
rect 144 2960 148 2962
rect 144 2954 148 2956
rect 144 2948 148 2950
rect 144 2942 148 2944
rect 144 2936 148 2938
rect 144 2930 148 2932
rect 144 2924 148 2926
rect 144 2918 148 2920
rect 144 2912 148 2914
rect 144 2906 148 2908
rect 144 2900 148 2902
rect 144 2894 148 2896
rect 144 2888 148 2890
rect 144 2882 148 2884
rect 144 2876 148 2878
rect 144 2870 148 2872
rect 144 2864 148 2866
rect 144 2858 148 2860
rect 144 2852 148 2854
rect 144 2846 148 2848
rect 148 2842 150 2846
rect 154 2842 156 2846
rect 160 2842 162 2846
rect 166 2842 168 2846
rect 172 2842 174 2846
rect 178 2842 180 2846
rect 184 2842 186 2846
rect 190 2842 192 2846
rect 196 2842 198 2846
rect 202 2842 204 2846
rect 208 2842 210 2846
rect 214 2842 216 2846
rect 220 2842 222 2846
rect 226 2842 228 2846
rect 232 2842 234 2846
rect 238 2842 240 2846
rect 244 2842 246 2846
rect 250 2842 252 2846
rect 256 2842 258 2846
rect 262 2842 264 2846
rect 268 2842 270 2846
rect 274 2842 276 2846
rect 280 2842 282 2846
rect 286 2842 288 2846
rect 292 2842 294 2846
rect 298 2842 300 2846
rect 304 2842 306 2846
rect 310 2842 312 2846
rect 316 2842 318 2846
rect 322 2842 324 2846
rect 328 2842 330 2846
rect 334 2842 336 2846
rect 340 2842 342 2846
rect 346 2842 348 2846
rect 352 2842 354 2846
rect 358 2842 360 2846
rect 364 2842 366 2846
rect 370 2842 372 2846
rect 376 2842 378 2846
rect 382 2842 384 2846
rect 388 2842 390 2846
rect 394 2842 396 2846
rect 400 2842 402 2846
rect 406 2842 408 2846
rect 412 2842 414 2846
rect 418 2842 420 2846
rect 424 2842 426 2846
rect 430 2842 432 2846
rect 436 2842 438 2846
rect 442 2842 444 2846
rect 448 2842 450 2846
rect 454 2842 456 2846
rect 460 2842 462 2846
rect 466 2842 468 2846
rect 472 2842 474 2846
rect 478 2842 480 2846
rect 484 2842 486 2846
rect 490 2842 492 2846
rect 496 2842 498 2846
rect 502 2842 504 2846
rect 508 2842 510 2846
rect 144 2840 148 2842
rect 144 2834 148 2836
rect 144 2828 148 2830
rect 144 2822 148 2824
rect 144 2816 148 2818
rect 144 2810 148 2812
rect 144 2804 148 2806
rect 144 2798 148 2800
rect 144 2792 148 2794
rect 144 2786 148 2788
rect 144 2780 148 2782
rect 144 2774 148 2776
rect 144 2768 148 2770
rect 144 2762 148 2764
rect 144 2756 148 2758
rect 144 2750 148 2752
rect 144 2744 148 2746
rect 144 2738 148 2740
rect 144 2732 148 2734
rect 144 2726 148 2728
rect 144 2720 148 2722
rect 4 2712 8 2716
rect 12 2712 63 2716
rect 72 2712 74 2716
rect 78 2712 80 2716
rect 84 2712 86 2716
rect 90 2712 92 2716
rect 101 2712 137 2716
rect 141 2714 148 2716
rect 141 2712 144 2714
rect 0 2710 144 2712
rect 4 2706 8 2710
rect 12 2706 63 2710
rect 72 2706 74 2710
rect 78 2706 80 2710
rect 84 2706 86 2710
rect 90 2706 92 2710
rect 101 2706 137 2710
rect 141 2708 148 2710
rect 141 2706 144 2708
rect 0 2704 144 2706
rect 4 2700 8 2704
rect 12 2700 63 2704
rect 72 2700 74 2704
rect 78 2700 80 2704
rect 84 2700 86 2704
rect 90 2700 92 2704
rect 101 2700 137 2704
rect 141 2702 148 2704
rect 141 2700 144 2702
rect 0 2698 144 2700
rect 4 2694 8 2698
rect 12 2694 63 2698
rect 72 2694 74 2698
rect 78 2694 80 2698
rect 84 2694 86 2698
rect 90 2694 92 2698
rect 101 2694 137 2698
rect 141 2696 148 2698
rect 141 2694 144 2696
rect 0 2692 144 2694
rect 4 2688 8 2692
rect 12 2688 63 2692
rect 72 2688 74 2692
rect 78 2688 80 2692
rect 84 2688 86 2692
rect 90 2688 92 2692
rect 101 2688 137 2692
rect 141 2690 148 2692
rect 141 2688 144 2690
rect 0 2686 144 2688
rect 4 2682 8 2686
rect 12 2682 63 2686
rect 72 2682 74 2686
rect 78 2682 80 2686
rect 84 2682 86 2686
rect 90 2682 92 2686
rect 101 2682 137 2686
rect 141 2684 148 2686
rect 141 2682 144 2684
rect 0 2680 144 2682
rect 4 2676 8 2680
rect 12 2676 63 2680
rect 72 2676 74 2680
rect 78 2676 80 2680
rect 84 2676 86 2680
rect 90 2676 92 2680
rect 101 2676 137 2680
rect 141 2678 148 2680
rect 141 2676 144 2678
rect 144 2672 148 2674
rect 4 2668 20 2672
rect 24 2668 26 2672
rect 30 2668 32 2672
rect 36 2668 38 2672
rect 42 2668 44 2672
rect 48 2671 100 2672
rect 48 2668 64 2671
rect 0 2667 64 2668
rect 68 2667 70 2671
rect 74 2667 76 2671
rect 80 2667 82 2671
rect 86 2667 89 2671
rect 93 2667 95 2671
rect 99 2667 100 2671
rect 0 2666 100 2667
rect 4 2662 14 2666
rect 18 2662 20 2666
rect 24 2662 26 2666
rect 30 2662 32 2666
rect 36 2662 38 2666
rect 42 2662 44 2666
rect 48 2665 100 2666
rect 48 2662 64 2665
rect 0 2661 64 2662
rect 68 2661 70 2665
rect 74 2661 76 2665
rect 80 2661 82 2665
rect 86 2661 89 2665
rect 93 2661 95 2665
rect 99 2661 100 2665
rect 0 2660 100 2661
rect 4 2656 14 2660
rect 18 2656 20 2660
rect 24 2656 26 2660
rect 30 2656 32 2660
rect 36 2656 38 2660
rect 42 2656 44 2660
rect 48 2659 100 2660
rect 48 2656 64 2659
rect 0 2655 64 2656
rect 68 2655 70 2659
rect 74 2655 76 2659
rect 80 2655 82 2659
rect 86 2655 89 2659
rect 93 2655 95 2659
rect 99 2655 100 2659
rect 0 2654 100 2655
rect 4 2650 14 2654
rect 18 2650 20 2654
rect 24 2650 26 2654
rect 30 2650 32 2654
rect 36 2650 38 2654
rect 42 2650 44 2654
rect 48 2653 100 2654
rect 48 2650 64 2653
rect 0 2649 64 2650
rect 68 2649 70 2653
rect 74 2649 76 2653
rect 80 2649 82 2653
rect 86 2649 89 2653
rect 93 2649 95 2653
rect 99 2649 100 2653
rect 0 2648 100 2649
rect 4 2644 14 2648
rect 18 2644 20 2648
rect 24 2644 26 2648
rect 30 2644 32 2648
rect 36 2644 38 2648
rect 42 2644 44 2648
rect 48 2647 100 2648
rect 48 2644 64 2647
rect 0 2643 64 2644
rect 68 2643 70 2647
rect 74 2643 76 2647
rect 80 2643 82 2647
rect 86 2643 89 2647
rect 93 2643 95 2647
rect 99 2643 100 2647
rect 0 2642 100 2643
rect 111 2668 112 2672
rect 116 2668 119 2672
rect 123 2668 125 2672
rect 107 2666 129 2668
rect 144 2666 148 2668
rect 111 2662 112 2666
rect 116 2662 119 2666
rect 123 2662 125 2666
rect 129 2662 131 2666
rect 107 2660 135 2662
rect 111 2656 112 2660
rect 116 2656 119 2660
rect 123 2656 125 2660
rect 129 2656 131 2660
rect 107 2654 135 2656
rect 111 2650 112 2654
rect 116 2650 119 2654
rect 123 2650 125 2654
rect 129 2650 131 2654
rect 107 2648 135 2650
rect 111 2644 112 2648
rect 116 2644 119 2648
rect 123 2644 125 2648
rect 129 2644 131 2648
rect 107 2642 135 2644
rect 4 2638 14 2642
rect 18 2638 20 2642
rect 24 2638 26 2642
rect 30 2638 32 2642
rect 36 2638 38 2642
rect 42 2638 44 2642
rect 111 2638 112 2642
rect 116 2638 119 2642
rect 123 2638 125 2642
rect 129 2638 131 2642
rect 0 2636 48 2638
rect 4 2632 14 2636
rect 18 2632 20 2636
rect 24 2632 26 2636
rect 30 2632 32 2636
rect 36 2632 38 2636
rect 42 2632 44 2636
rect 52 2634 53 2638
rect 57 2634 58 2638
rect 52 2633 58 2634
rect 52 2629 53 2633
rect 57 2629 58 2633
rect 107 2636 135 2638
rect 111 2632 112 2636
rect 116 2632 119 2636
rect 123 2632 125 2636
rect 129 2632 131 2636
rect 144 2660 148 2662
rect 144 2654 148 2656
rect 144 2648 148 2650
rect 144 2642 148 2644
rect 144 2636 148 2638
rect 52 2628 58 2629
rect 4 2624 53 2628
rect 57 2624 58 2628
rect 4 2623 58 2624
rect 4 2619 53 2623
rect 57 2619 58 2623
rect 144 2630 148 2632
rect 144 2624 148 2626
rect 4 2591 53 2595
rect 57 2591 58 2595
rect 4 2590 58 2591
rect 4 2586 53 2590
rect 57 2586 58 2590
rect 52 2585 58 2586
rect 4 2578 14 2582
rect 18 2578 20 2582
rect 24 2578 26 2582
rect 30 2578 32 2582
rect 36 2578 38 2582
rect 42 2578 44 2582
rect 0 2576 48 2578
rect 52 2581 53 2585
rect 57 2581 58 2585
rect 144 2588 148 2590
rect 144 2582 148 2584
rect 52 2580 58 2581
rect 52 2576 53 2580
rect 57 2576 58 2580
rect 111 2578 112 2582
rect 116 2578 119 2582
rect 123 2578 125 2582
rect 129 2578 131 2582
rect 107 2576 135 2578
rect 4 2572 14 2576
rect 18 2572 20 2576
rect 24 2572 26 2576
rect 30 2572 32 2576
rect 36 2572 38 2576
rect 42 2572 44 2576
rect 111 2572 112 2576
rect 116 2572 119 2576
rect 123 2572 125 2576
rect 129 2572 131 2576
rect 0 2571 100 2572
rect 0 2570 64 2571
rect 4 2566 14 2570
rect 18 2566 20 2570
rect 24 2566 26 2570
rect 30 2566 32 2570
rect 36 2566 38 2570
rect 42 2566 44 2570
rect 48 2567 64 2570
rect 68 2567 70 2571
rect 74 2567 76 2571
rect 80 2567 82 2571
rect 86 2567 89 2571
rect 93 2567 95 2571
rect 99 2567 100 2571
rect 48 2566 100 2567
rect 0 2565 100 2566
rect 0 2564 64 2565
rect 4 2560 14 2564
rect 18 2560 20 2564
rect 24 2560 26 2564
rect 30 2560 32 2564
rect 36 2560 38 2564
rect 42 2560 44 2564
rect 48 2561 64 2564
rect 68 2561 70 2565
rect 74 2561 76 2565
rect 80 2561 82 2565
rect 86 2561 89 2565
rect 93 2561 95 2565
rect 99 2561 100 2565
rect 48 2560 100 2561
rect 0 2559 100 2560
rect 0 2558 64 2559
rect 4 2554 14 2558
rect 18 2554 20 2558
rect 24 2554 26 2558
rect 30 2554 32 2558
rect 36 2554 38 2558
rect 42 2554 44 2558
rect 48 2555 64 2558
rect 68 2555 70 2559
rect 74 2555 76 2559
rect 80 2555 82 2559
rect 86 2555 89 2559
rect 93 2555 95 2559
rect 99 2555 100 2559
rect 48 2554 100 2555
rect 0 2553 100 2554
rect 0 2552 64 2553
rect 4 2548 14 2552
rect 18 2548 20 2552
rect 24 2548 26 2552
rect 30 2548 32 2552
rect 36 2548 38 2552
rect 42 2548 44 2552
rect 48 2549 64 2552
rect 68 2549 70 2553
rect 74 2549 76 2553
rect 80 2549 82 2553
rect 86 2549 89 2553
rect 93 2549 95 2553
rect 99 2549 100 2553
rect 48 2548 100 2549
rect 0 2547 100 2548
rect 0 2546 64 2547
rect 4 2542 20 2546
rect 24 2542 26 2546
rect 30 2542 32 2546
rect 36 2542 38 2546
rect 42 2542 44 2546
rect 48 2543 64 2546
rect 68 2543 70 2547
rect 74 2543 76 2547
rect 80 2543 82 2547
rect 86 2543 89 2547
rect 93 2543 95 2547
rect 99 2543 100 2547
rect 48 2542 100 2543
rect 107 2570 135 2572
rect 111 2566 112 2570
rect 116 2566 119 2570
rect 123 2566 125 2570
rect 129 2566 131 2570
rect 107 2564 135 2566
rect 111 2560 112 2564
rect 116 2560 119 2564
rect 123 2560 125 2564
rect 129 2560 131 2564
rect 107 2558 135 2560
rect 111 2554 112 2558
rect 116 2554 119 2558
rect 123 2554 125 2558
rect 129 2554 131 2558
rect 107 2552 135 2554
rect 111 2548 112 2552
rect 116 2548 119 2552
rect 123 2548 125 2552
rect 129 2548 131 2552
rect 144 2576 148 2578
rect 144 2570 148 2572
rect 144 2564 148 2566
rect 144 2558 148 2560
rect 144 2552 148 2554
rect 107 2546 129 2548
rect 111 2542 112 2546
rect 116 2542 119 2546
rect 123 2542 125 2546
rect 144 2546 148 2548
rect 144 2540 148 2542
rect 4 2534 8 2538
rect 12 2534 63 2538
rect 72 2534 74 2538
rect 78 2534 80 2538
rect 84 2534 86 2538
rect 90 2534 92 2538
rect 101 2534 137 2538
rect 141 2536 144 2538
rect 141 2534 148 2536
rect 0 2532 144 2534
rect 4 2528 8 2532
rect 12 2528 63 2532
rect 72 2528 74 2532
rect 78 2528 80 2532
rect 84 2528 86 2532
rect 90 2528 92 2532
rect 101 2528 137 2532
rect 141 2530 144 2532
rect 141 2528 148 2530
rect 0 2526 144 2528
rect 4 2522 8 2526
rect 12 2522 63 2526
rect 72 2522 74 2526
rect 78 2522 80 2526
rect 84 2522 86 2526
rect 90 2522 92 2526
rect 101 2522 137 2526
rect 141 2524 144 2526
rect 141 2522 148 2524
rect 0 2520 144 2522
rect 4 2516 8 2520
rect 12 2516 63 2520
rect 72 2516 74 2520
rect 78 2516 80 2520
rect 84 2516 86 2520
rect 90 2516 92 2520
rect 101 2516 137 2520
rect 141 2518 144 2520
rect 141 2516 148 2518
rect 0 2514 144 2516
rect 4 2510 8 2514
rect 12 2510 63 2514
rect 72 2510 74 2514
rect 78 2510 80 2514
rect 84 2510 86 2514
rect 90 2510 92 2514
rect 101 2510 137 2514
rect 141 2512 144 2514
rect 141 2510 148 2512
rect 0 2508 144 2510
rect 4 2504 8 2508
rect 12 2504 63 2508
rect 72 2504 74 2508
rect 78 2504 80 2508
rect 84 2504 86 2508
rect 90 2504 92 2508
rect 101 2504 137 2508
rect 141 2506 144 2508
rect 141 2504 148 2506
rect 0 2502 144 2504
rect 4 2498 8 2502
rect 12 2498 63 2502
rect 72 2498 74 2502
rect 78 2498 80 2502
rect 84 2498 86 2502
rect 90 2498 92 2502
rect 101 2498 137 2502
rect 141 2500 144 2502
rect 141 2498 148 2500
rect 144 2492 148 2494
rect 144 2486 148 2488
rect 144 2480 148 2482
rect 144 2474 148 2476
rect 144 2468 148 2470
rect 144 2462 148 2464
rect 144 2456 148 2458
rect 144 2450 148 2452
rect 144 2444 148 2446
rect 144 2438 148 2440
rect 144 2432 148 2434
rect 144 2426 148 2428
rect 144 2420 148 2422
rect 144 2414 148 2416
rect 144 2408 148 2410
rect 144 2402 148 2404
rect 144 2396 148 2398
rect 144 2390 148 2392
rect 144 2384 148 2386
rect 144 2378 148 2380
rect 144 2372 148 2374
rect 148 2368 150 2372
rect 154 2368 156 2372
rect 160 2368 162 2372
rect 166 2368 168 2372
rect 172 2368 174 2372
rect 178 2368 180 2372
rect 184 2368 186 2372
rect 190 2368 192 2372
rect 196 2368 198 2372
rect 202 2368 204 2372
rect 208 2368 210 2372
rect 214 2368 216 2372
rect 220 2368 222 2372
rect 226 2368 228 2372
rect 232 2368 234 2372
rect 238 2368 240 2372
rect 244 2368 246 2372
rect 250 2368 252 2372
rect 256 2368 258 2372
rect 262 2368 264 2372
rect 268 2368 270 2372
rect 274 2368 276 2372
rect 280 2368 282 2372
rect 286 2368 288 2372
rect 292 2368 294 2372
rect 298 2368 300 2372
rect 304 2368 306 2372
rect 310 2368 312 2372
rect 316 2368 318 2372
rect 322 2368 324 2372
rect 328 2368 330 2372
rect 334 2368 336 2372
rect 340 2368 342 2372
rect 346 2368 348 2372
rect 352 2368 354 2372
rect 358 2368 360 2372
rect 364 2368 366 2372
rect 370 2368 372 2372
rect 376 2368 378 2372
rect 382 2368 384 2372
rect 388 2368 390 2372
rect 394 2368 396 2372
rect 400 2368 402 2372
rect 406 2368 408 2372
rect 412 2368 414 2372
rect 418 2368 420 2372
rect 424 2368 426 2372
rect 430 2368 432 2372
rect 436 2368 438 2372
rect 442 2368 444 2372
rect 448 2368 450 2372
rect 454 2368 456 2372
rect 460 2368 462 2372
rect 466 2368 468 2372
rect 472 2368 474 2372
rect 478 2368 480 2372
rect 484 2368 486 2372
rect 490 2368 492 2372
rect 496 2368 498 2372
rect 502 2368 504 2372
rect 508 2368 510 2372
rect 144 2366 148 2368
rect 144 2360 148 2362
rect 144 2354 148 2356
rect 144 2348 148 2350
rect 144 2342 148 2344
rect 144 2336 148 2338
rect 144 2330 148 2332
rect 144 2324 148 2326
rect 144 2318 148 2320
rect 144 2312 148 2314
rect 144 2306 148 2308
rect 144 2300 148 2302
rect 144 2294 148 2296
rect 144 2288 148 2290
rect 144 2282 148 2284
rect 144 2276 148 2278
rect 144 2270 148 2272
rect 144 2264 148 2266
rect 144 2258 148 2260
rect 144 2252 148 2254
rect 144 2246 148 2248
rect 4 2238 8 2242
rect 12 2238 63 2242
rect 72 2238 74 2242
rect 78 2238 80 2242
rect 84 2238 86 2242
rect 90 2238 92 2242
rect 101 2238 137 2242
rect 141 2240 148 2242
rect 141 2238 144 2240
rect 0 2236 144 2238
rect 4 2232 8 2236
rect 12 2232 63 2236
rect 72 2232 74 2236
rect 78 2232 80 2236
rect 84 2232 86 2236
rect 90 2232 92 2236
rect 101 2232 137 2236
rect 141 2234 148 2236
rect 141 2232 144 2234
rect 0 2230 144 2232
rect 4 2226 8 2230
rect 12 2226 63 2230
rect 72 2226 74 2230
rect 78 2226 80 2230
rect 84 2226 86 2230
rect 90 2226 92 2230
rect 101 2226 137 2230
rect 141 2228 148 2230
rect 141 2226 144 2228
rect 0 2224 144 2226
rect 4 2220 8 2224
rect 12 2220 63 2224
rect 72 2220 74 2224
rect 78 2220 80 2224
rect 84 2220 86 2224
rect 90 2220 92 2224
rect 101 2220 137 2224
rect 141 2222 148 2224
rect 141 2220 144 2222
rect 0 2218 144 2220
rect 4 2214 8 2218
rect 12 2214 63 2218
rect 72 2214 74 2218
rect 78 2214 80 2218
rect 84 2214 86 2218
rect 90 2214 92 2218
rect 101 2214 137 2218
rect 141 2216 148 2218
rect 141 2214 144 2216
rect 0 2212 144 2214
rect 4 2208 8 2212
rect 12 2208 63 2212
rect 72 2208 74 2212
rect 78 2208 80 2212
rect 84 2208 86 2212
rect 90 2208 92 2212
rect 101 2208 137 2212
rect 141 2210 148 2212
rect 141 2208 144 2210
rect 0 2206 144 2208
rect 4 2202 8 2206
rect 12 2202 63 2206
rect 72 2202 74 2206
rect 78 2202 80 2206
rect 84 2202 86 2206
rect 90 2202 92 2206
rect 101 2202 137 2206
rect 141 2204 148 2206
rect 141 2202 144 2204
rect 144 2198 148 2200
rect 4 2194 20 2198
rect 24 2194 26 2198
rect 30 2194 32 2198
rect 36 2194 38 2198
rect 42 2194 44 2198
rect 48 2197 100 2198
rect 48 2194 64 2197
rect 0 2193 64 2194
rect 68 2193 70 2197
rect 74 2193 76 2197
rect 80 2193 82 2197
rect 86 2193 89 2197
rect 93 2193 95 2197
rect 99 2193 100 2197
rect 0 2192 100 2193
rect 4 2188 14 2192
rect 18 2188 20 2192
rect 24 2188 26 2192
rect 30 2188 32 2192
rect 36 2188 38 2192
rect 42 2188 44 2192
rect 48 2191 100 2192
rect 48 2188 64 2191
rect 0 2187 64 2188
rect 68 2187 70 2191
rect 74 2187 76 2191
rect 80 2187 82 2191
rect 86 2187 89 2191
rect 93 2187 95 2191
rect 99 2187 100 2191
rect 0 2186 100 2187
rect 4 2182 14 2186
rect 18 2182 20 2186
rect 24 2182 26 2186
rect 30 2182 32 2186
rect 36 2182 38 2186
rect 42 2182 44 2186
rect 48 2185 100 2186
rect 48 2182 64 2185
rect 0 2181 64 2182
rect 68 2181 70 2185
rect 74 2181 76 2185
rect 80 2181 82 2185
rect 86 2181 89 2185
rect 93 2181 95 2185
rect 99 2181 100 2185
rect 0 2180 100 2181
rect 4 2176 14 2180
rect 18 2176 20 2180
rect 24 2176 26 2180
rect 30 2176 32 2180
rect 36 2176 38 2180
rect 42 2176 44 2180
rect 48 2179 100 2180
rect 48 2176 64 2179
rect 0 2175 64 2176
rect 68 2175 70 2179
rect 74 2175 76 2179
rect 80 2175 82 2179
rect 86 2175 89 2179
rect 93 2175 95 2179
rect 99 2175 100 2179
rect 0 2174 100 2175
rect 4 2170 14 2174
rect 18 2170 20 2174
rect 24 2170 26 2174
rect 30 2170 32 2174
rect 36 2170 38 2174
rect 42 2170 44 2174
rect 48 2173 100 2174
rect 48 2170 64 2173
rect 0 2169 64 2170
rect 68 2169 70 2173
rect 74 2169 76 2173
rect 80 2169 82 2173
rect 86 2169 89 2173
rect 93 2169 95 2173
rect 99 2169 100 2173
rect 0 2168 100 2169
rect 111 2194 112 2198
rect 116 2194 119 2198
rect 123 2194 125 2198
rect 107 2192 129 2194
rect 144 2192 148 2194
rect 111 2188 112 2192
rect 116 2188 119 2192
rect 123 2188 125 2192
rect 129 2188 131 2192
rect 107 2186 135 2188
rect 111 2182 112 2186
rect 116 2182 119 2186
rect 123 2182 125 2186
rect 129 2182 131 2186
rect 107 2180 135 2182
rect 111 2176 112 2180
rect 116 2176 119 2180
rect 123 2176 125 2180
rect 129 2176 131 2180
rect 107 2174 135 2176
rect 111 2170 112 2174
rect 116 2170 119 2174
rect 123 2170 125 2174
rect 129 2170 131 2174
rect 107 2168 135 2170
rect 4 2164 14 2168
rect 18 2164 20 2168
rect 24 2164 26 2168
rect 30 2164 32 2168
rect 36 2164 38 2168
rect 42 2164 44 2168
rect 111 2164 112 2168
rect 116 2164 119 2168
rect 123 2164 125 2168
rect 129 2164 131 2168
rect 0 2162 48 2164
rect 4 2158 14 2162
rect 18 2158 20 2162
rect 24 2158 26 2162
rect 30 2158 32 2162
rect 36 2158 38 2162
rect 42 2158 44 2162
rect 52 2160 53 2164
rect 57 2160 58 2164
rect 52 2159 58 2160
rect 52 2155 53 2159
rect 57 2155 58 2159
rect 107 2162 135 2164
rect 111 2158 112 2162
rect 116 2158 119 2162
rect 123 2158 125 2162
rect 129 2158 131 2162
rect 144 2186 148 2188
rect 144 2180 148 2182
rect 144 2174 148 2176
rect 144 2168 148 2170
rect 144 2162 148 2164
rect 52 2154 58 2155
rect 4 2150 53 2154
rect 57 2150 58 2154
rect 4 2149 58 2150
rect 4 2145 53 2149
rect 57 2145 58 2149
rect 144 2156 148 2158
rect 144 2150 148 2152
rect 4 2117 53 2121
rect 57 2117 58 2121
rect 4 2116 58 2117
rect 4 2112 53 2116
rect 57 2112 58 2116
rect 52 2111 58 2112
rect 4 2104 14 2108
rect 18 2104 20 2108
rect 24 2104 26 2108
rect 30 2104 32 2108
rect 36 2104 38 2108
rect 42 2104 44 2108
rect 0 2102 48 2104
rect 52 2107 53 2111
rect 57 2107 58 2111
rect 144 2114 148 2116
rect 144 2108 148 2110
rect 52 2106 58 2107
rect 52 2102 53 2106
rect 57 2102 58 2106
rect 111 2104 112 2108
rect 116 2104 119 2108
rect 123 2104 125 2108
rect 129 2104 131 2108
rect 107 2102 135 2104
rect 4 2098 14 2102
rect 18 2098 20 2102
rect 24 2098 26 2102
rect 30 2098 32 2102
rect 36 2098 38 2102
rect 42 2098 44 2102
rect 111 2098 112 2102
rect 116 2098 119 2102
rect 123 2098 125 2102
rect 129 2098 131 2102
rect 0 2097 100 2098
rect 0 2096 64 2097
rect 4 2092 14 2096
rect 18 2092 20 2096
rect 24 2092 26 2096
rect 30 2092 32 2096
rect 36 2092 38 2096
rect 42 2092 44 2096
rect 48 2093 64 2096
rect 68 2093 70 2097
rect 74 2093 76 2097
rect 80 2093 82 2097
rect 86 2093 89 2097
rect 93 2093 95 2097
rect 99 2093 100 2097
rect 48 2092 100 2093
rect 0 2091 100 2092
rect 0 2090 64 2091
rect 4 2086 14 2090
rect 18 2086 20 2090
rect 24 2086 26 2090
rect 30 2086 32 2090
rect 36 2086 38 2090
rect 42 2086 44 2090
rect 48 2087 64 2090
rect 68 2087 70 2091
rect 74 2087 76 2091
rect 80 2087 82 2091
rect 86 2087 89 2091
rect 93 2087 95 2091
rect 99 2087 100 2091
rect 48 2086 100 2087
rect 0 2085 100 2086
rect 0 2084 64 2085
rect 4 2080 14 2084
rect 18 2080 20 2084
rect 24 2080 26 2084
rect 30 2080 32 2084
rect 36 2080 38 2084
rect 42 2080 44 2084
rect 48 2081 64 2084
rect 68 2081 70 2085
rect 74 2081 76 2085
rect 80 2081 82 2085
rect 86 2081 89 2085
rect 93 2081 95 2085
rect 99 2081 100 2085
rect 48 2080 100 2081
rect 0 2079 100 2080
rect 0 2078 64 2079
rect 4 2074 14 2078
rect 18 2074 20 2078
rect 24 2074 26 2078
rect 30 2074 32 2078
rect 36 2074 38 2078
rect 42 2074 44 2078
rect 48 2075 64 2078
rect 68 2075 70 2079
rect 74 2075 76 2079
rect 80 2075 82 2079
rect 86 2075 89 2079
rect 93 2075 95 2079
rect 99 2075 100 2079
rect 48 2074 100 2075
rect 0 2073 100 2074
rect 0 2072 64 2073
rect 4 2068 20 2072
rect 24 2068 26 2072
rect 30 2068 32 2072
rect 36 2068 38 2072
rect 42 2068 44 2072
rect 48 2069 64 2072
rect 68 2069 70 2073
rect 74 2069 76 2073
rect 80 2069 82 2073
rect 86 2069 89 2073
rect 93 2069 95 2073
rect 99 2069 100 2073
rect 48 2068 100 2069
rect 107 2096 135 2098
rect 111 2092 112 2096
rect 116 2092 119 2096
rect 123 2092 125 2096
rect 129 2092 131 2096
rect 107 2090 135 2092
rect 111 2086 112 2090
rect 116 2086 119 2090
rect 123 2086 125 2090
rect 129 2086 131 2090
rect 107 2084 135 2086
rect 111 2080 112 2084
rect 116 2080 119 2084
rect 123 2080 125 2084
rect 129 2080 131 2084
rect 107 2078 135 2080
rect 111 2074 112 2078
rect 116 2074 119 2078
rect 123 2074 125 2078
rect 129 2074 131 2078
rect 144 2102 148 2104
rect 144 2096 148 2098
rect 144 2090 148 2092
rect 144 2084 148 2086
rect 144 2078 148 2080
rect 107 2072 129 2074
rect 111 2068 112 2072
rect 116 2068 119 2072
rect 123 2068 125 2072
rect 144 2072 148 2074
rect 144 2066 148 2068
rect 4 2060 8 2064
rect 12 2060 63 2064
rect 72 2060 74 2064
rect 78 2060 80 2064
rect 84 2060 86 2064
rect 90 2060 92 2064
rect 101 2060 137 2064
rect 141 2062 144 2064
rect 141 2060 148 2062
rect 0 2058 144 2060
rect 4 2054 8 2058
rect 12 2054 63 2058
rect 72 2054 74 2058
rect 78 2054 80 2058
rect 84 2054 86 2058
rect 90 2054 92 2058
rect 101 2054 137 2058
rect 141 2056 144 2058
rect 141 2054 148 2056
rect 0 2052 144 2054
rect 4 2048 8 2052
rect 12 2048 63 2052
rect 72 2048 74 2052
rect 78 2048 80 2052
rect 84 2048 86 2052
rect 90 2048 92 2052
rect 101 2048 137 2052
rect 141 2050 144 2052
rect 141 2048 148 2050
rect 0 2046 144 2048
rect 4 2042 8 2046
rect 12 2042 63 2046
rect 72 2042 74 2046
rect 78 2042 80 2046
rect 84 2042 86 2046
rect 90 2042 92 2046
rect 101 2042 137 2046
rect 141 2044 144 2046
rect 141 2042 148 2044
rect 0 2040 144 2042
rect 4 2036 8 2040
rect 12 2036 63 2040
rect 72 2036 74 2040
rect 78 2036 80 2040
rect 84 2036 86 2040
rect 90 2036 92 2040
rect 101 2036 137 2040
rect 141 2038 144 2040
rect 141 2036 148 2038
rect 0 2034 144 2036
rect 4 2030 8 2034
rect 12 2030 63 2034
rect 72 2030 74 2034
rect 78 2030 80 2034
rect 84 2030 86 2034
rect 90 2030 92 2034
rect 101 2030 137 2034
rect 141 2032 144 2034
rect 141 2030 148 2032
rect 0 2028 144 2030
rect 4 2024 8 2028
rect 12 2024 63 2028
rect 72 2024 74 2028
rect 78 2024 80 2028
rect 84 2024 86 2028
rect 90 2024 92 2028
rect 101 2024 137 2028
rect 141 2026 144 2028
rect 141 2024 148 2026
rect 144 2018 148 2020
rect 144 2012 148 2014
rect 144 2006 148 2008
rect 144 2000 148 2002
rect 144 1994 148 1996
rect 144 1988 148 1990
rect 144 1982 148 1984
rect 144 1976 148 1978
rect 144 1970 148 1972
rect 144 1964 148 1966
rect 144 1958 148 1960
rect 144 1952 148 1954
rect 144 1946 148 1948
rect 144 1940 148 1942
rect 144 1934 148 1936
rect 144 1928 148 1930
rect 144 1922 148 1924
rect 144 1916 148 1918
rect 144 1910 148 1912
rect 144 1904 148 1906
rect 144 1898 148 1900
rect 148 1894 150 1898
rect 154 1894 156 1898
rect 160 1894 162 1898
rect 166 1894 168 1898
rect 172 1894 174 1898
rect 178 1894 180 1898
rect 184 1894 186 1898
rect 190 1894 192 1898
rect 196 1894 198 1898
rect 202 1894 204 1898
rect 208 1894 210 1898
rect 214 1894 216 1898
rect 220 1894 222 1898
rect 226 1894 228 1898
rect 232 1894 234 1898
rect 238 1894 240 1898
rect 244 1894 246 1898
rect 250 1894 252 1898
rect 256 1894 258 1898
rect 262 1894 264 1898
rect 268 1894 270 1898
rect 274 1894 276 1898
rect 280 1894 282 1898
rect 286 1894 288 1898
rect 292 1894 294 1898
rect 298 1894 300 1898
rect 304 1894 306 1898
rect 310 1894 312 1898
rect 316 1894 318 1898
rect 322 1894 324 1898
rect 328 1894 330 1898
rect 334 1894 336 1898
rect 340 1894 342 1898
rect 346 1894 348 1898
rect 352 1894 354 1898
rect 358 1894 360 1898
rect 364 1894 366 1898
rect 370 1894 372 1898
rect 376 1894 378 1898
rect 382 1894 384 1898
rect 388 1894 390 1898
rect 394 1894 396 1898
rect 400 1894 402 1898
rect 406 1894 408 1898
rect 412 1894 414 1898
rect 418 1894 420 1898
rect 424 1894 426 1898
rect 430 1894 432 1898
rect 436 1894 438 1898
rect 442 1894 444 1898
rect 448 1894 450 1898
rect 454 1894 456 1898
rect 460 1894 462 1898
rect 466 1894 468 1898
rect 472 1894 474 1898
rect 478 1894 480 1898
rect 484 1894 486 1898
rect 490 1894 492 1898
rect 496 1894 498 1898
rect 502 1894 504 1898
rect 508 1894 510 1898
rect 144 1892 148 1894
rect 144 1886 148 1888
rect 144 1880 148 1882
rect 144 1874 148 1876
rect 144 1868 148 1870
rect 144 1862 148 1864
rect 144 1856 148 1858
rect 144 1850 148 1852
rect 144 1844 148 1846
rect 144 1838 148 1840
rect 144 1832 148 1834
rect 144 1826 148 1828
rect 144 1820 148 1822
rect 144 1814 148 1816
rect 144 1808 148 1810
rect 144 1802 148 1804
rect 144 1796 148 1798
rect 144 1790 148 1792
rect 144 1784 148 1786
rect 144 1778 148 1780
rect 144 1772 148 1774
rect 4 1764 8 1768
rect 12 1764 63 1768
rect 72 1764 74 1768
rect 78 1764 80 1768
rect 84 1764 86 1768
rect 90 1764 92 1768
rect 101 1764 137 1768
rect 141 1766 148 1768
rect 141 1764 144 1766
rect 0 1762 144 1764
rect 4 1758 8 1762
rect 12 1758 63 1762
rect 72 1758 74 1762
rect 78 1758 80 1762
rect 84 1758 86 1762
rect 90 1758 92 1762
rect 101 1758 137 1762
rect 141 1760 148 1762
rect 141 1758 144 1760
rect 0 1756 144 1758
rect 4 1752 8 1756
rect 12 1752 63 1756
rect 72 1752 74 1756
rect 78 1752 80 1756
rect 84 1752 86 1756
rect 90 1752 92 1756
rect 101 1752 137 1756
rect 141 1754 148 1756
rect 141 1752 144 1754
rect 0 1750 144 1752
rect 4 1746 8 1750
rect 12 1746 63 1750
rect 72 1746 74 1750
rect 78 1746 80 1750
rect 84 1746 86 1750
rect 90 1746 92 1750
rect 101 1746 137 1750
rect 141 1748 148 1750
rect 141 1746 144 1748
rect 0 1744 144 1746
rect 4 1740 8 1744
rect 12 1740 63 1744
rect 72 1740 74 1744
rect 78 1740 80 1744
rect 84 1740 86 1744
rect 90 1740 92 1744
rect 101 1740 137 1744
rect 141 1742 148 1744
rect 141 1740 144 1742
rect 0 1738 144 1740
rect 4 1734 8 1738
rect 12 1734 63 1738
rect 72 1734 74 1738
rect 78 1734 80 1738
rect 84 1734 86 1738
rect 90 1734 92 1738
rect 101 1734 137 1738
rect 141 1736 148 1738
rect 141 1734 144 1736
rect 0 1732 144 1734
rect 4 1728 8 1732
rect 12 1728 63 1732
rect 72 1728 74 1732
rect 78 1728 80 1732
rect 84 1728 86 1732
rect 90 1728 92 1732
rect 101 1728 137 1732
rect 141 1730 148 1732
rect 141 1728 144 1730
rect 144 1724 148 1726
rect 4 1720 20 1724
rect 24 1720 26 1724
rect 30 1720 32 1724
rect 36 1720 38 1724
rect 42 1720 44 1724
rect 48 1723 100 1724
rect 48 1720 64 1723
rect 0 1719 64 1720
rect 68 1719 70 1723
rect 74 1719 76 1723
rect 80 1719 82 1723
rect 86 1719 89 1723
rect 93 1719 95 1723
rect 99 1719 100 1723
rect 0 1718 100 1719
rect 4 1714 14 1718
rect 18 1714 20 1718
rect 24 1714 26 1718
rect 30 1714 32 1718
rect 36 1714 38 1718
rect 42 1714 44 1718
rect 48 1717 100 1718
rect 48 1714 64 1717
rect 0 1713 64 1714
rect 68 1713 70 1717
rect 74 1713 76 1717
rect 80 1713 82 1717
rect 86 1713 89 1717
rect 93 1713 95 1717
rect 99 1713 100 1717
rect 0 1712 100 1713
rect 4 1708 14 1712
rect 18 1708 20 1712
rect 24 1708 26 1712
rect 30 1708 32 1712
rect 36 1708 38 1712
rect 42 1708 44 1712
rect 48 1711 100 1712
rect 48 1708 64 1711
rect 0 1707 64 1708
rect 68 1707 70 1711
rect 74 1707 76 1711
rect 80 1707 82 1711
rect 86 1707 89 1711
rect 93 1707 95 1711
rect 99 1707 100 1711
rect 0 1706 100 1707
rect 4 1702 14 1706
rect 18 1702 20 1706
rect 24 1702 26 1706
rect 30 1702 32 1706
rect 36 1702 38 1706
rect 42 1702 44 1706
rect 48 1705 100 1706
rect 48 1702 64 1705
rect 0 1701 64 1702
rect 68 1701 70 1705
rect 74 1701 76 1705
rect 80 1701 82 1705
rect 86 1701 89 1705
rect 93 1701 95 1705
rect 99 1701 100 1705
rect 0 1700 100 1701
rect 4 1696 14 1700
rect 18 1696 20 1700
rect 24 1696 26 1700
rect 30 1696 32 1700
rect 36 1696 38 1700
rect 42 1696 44 1700
rect 48 1699 100 1700
rect 48 1696 64 1699
rect 0 1695 64 1696
rect 68 1695 70 1699
rect 74 1695 76 1699
rect 80 1695 82 1699
rect 86 1695 89 1699
rect 93 1695 95 1699
rect 99 1695 100 1699
rect 0 1694 100 1695
rect 111 1720 112 1724
rect 116 1720 119 1724
rect 123 1720 125 1724
rect 107 1718 129 1720
rect 144 1718 148 1720
rect 111 1714 112 1718
rect 116 1714 119 1718
rect 123 1714 125 1718
rect 129 1714 131 1718
rect 107 1712 135 1714
rect 111 1708 112 1712
rect 116 1708 119 1712
rect 123 1708 125 1712
rect 129 1708 131 1712
rect 107 1706 135 1708
rect 111 1702 112 1706
rect 116 1702 119 1706
rect 123 1702 125 1706
rect 129 1702 131 1706
rect 107 1700 135 1702
rect 111 1696 112 1700
rect 116 1696 119 1700
rect 123 1696 125 1700
rect 129 1696 131 1700
rect 107 1694 135 1696
rect 4 1690 14 1694
rect 18 1690 20 1694
rect 24 1690 26 1694
rect 30 1690 32 1694
rect 36 1690 38 1694
rect 42 1690 44 1694
rect 111 1690 112 1694
rect 116 1690 119 1694
rect 123 1690 125 1694
rect 129 1690 131 1694
rect 0 1688 48 1690
rect 4 1684 14 1688
rect 18 1684 20 1688
rect 24 1684 26 1688
rect 30 1684 32 1688
rect 36 1684 38 1688
rect 42 1684 44 1688
rect 52 1686 53 1690
rect 57 1686 58 1690
rect 52 1685 58 1686
rect 52 1681 53 1685
rect 57 1681 58 1685
rect 107 1688 135 1690
rect 111 1684 112 1688
rect 116 1684 119 1688
rect 123 1684 125 1688
rect 129 1684 131 1688
rect 144 1712 148 1714
rect 144 1706 148 1708
rect 144 1700 148 1702
rect 144 1694 148 1696
rect 144 1688 148 1690
rect 52 1680 58 1681
rect 4 1676 53 1680
rect 57 1676 58 1680
rect 4 1675 58 1676
rect 4 1671 53 1675
rect 57 1671 58 1675
rect 144 1682 148 1684
rect 144 1676 148 1678
rect 4 1643 53 1647
rect 57 1643 58 1647
rect 4 1642 58 1643
rect 4 1638 53 1642
rect 57 1638 58 1642
rect 52 1637 58 1638
rect 4 1630 14 1634
rect 18 1630 20 1634
rect 24 1630 26 1634
rect 30 1630 32 1634
rect 36 1630 38 1634
rect 42 1630 44 1634
rect 0 1628 48 1630
rect 52 1633 53 1637
rect 57 1633 58 1637
rect 144 1640 148 1642
rect 144 1634 148 1636
rect 52 1632 58 1633
rect 52 1628 53 1632
rect 57 1628 58 1632
rect 111 1630 112 1634
rect 116 1630 119 1634
rect 123 1630 125 1634
rect 129 1630 131 1634
rect 107 1628 135 1630
rect 4 1624 14 1628
rect 18 1624 20 1628
rect 24 1624 26 1628
rect 30 1624 32 1628
rect 36 1624 38 1628
rect 42 1624 44 1628
rect 111 1624 112 1628
rect 116 1624 119 1628
rect 123 1624 125 1628
rect 129 1624 131 1628
rect 0 1623 100 1624
rect 0 1622 64 1623
rect 4 1618 14 1622
rect 18 1618 20 1622
rect 24 1618 26 1622
rect 30 1618 32 1622
rect 36 1618 38 1622
rect 42 1618 44 1622
rect 48 1619 64 1622
rect 68 1619 70 1623
rect 74 1619 76 1623
rect 80 1619 82 1623
rect 86 1619 89 1623
rect 93 1619 95 1623
rect 99 1619 100 1623
rect 48 1618 100 1619
rect 0 1617 100 1618
rect 0 1616 64 1617
rect 4 1612 14 1616
rect 18 1612 20 1616
rect 24 1612 26 1616
rect 30 1612 32 1616
rect 36 1612 38 1616
rect 42 1612 44 1616
rect 48 1613 64 1616
rect 68 1613 70 1617
rect 74 1613 76 1617
rect 80 1613 82 1617
rect 86 1613 89 1617
rect 93 1613 95 1617
rect 99 1613 100 1617
rect 48 1612 100 1613
rect 0 1611 100 1612
rect 0 1610 64 1611
rect 4 1606 14 1610
rect 18 1606 20 1610
rect 24 1606 26 1610
rect 30 1606 32 1610
rect 36 1606 38 1610
rect 42 1606 44 1610
rect 48 1607 64 1610
rect 68 1607 70 1611
rect 74 1607 76 1611
rect 80 1607 82 1611
rect 86 1607 89 1611
rect 93 1607 95 1611
rect 99 1607 100 1611
rect 48 1606 100 1607
rect 0 1605 100 1606
rect 0 1604 64 1605
rect 4 1600 14 1604
rect 18 1600 20 1604
rect 24 1600 26 1604
rect 30 1600 32 1604
rect 36 1600 38 1604
rect 42 1600 44 1604
rect 48 1601 64 1604
rect 68 1601 70 1605
rect 74 1601 76 1605
rect 80 1601 82 1605
rect 86 1601 89 1605
rect 93 1601 95 1605
rect 99 1601 100 1605
rect 48 1600 100 1601
rect 0 1599 100 1600
rect 0 1598 64 1599
rect 4 1594 20 1598
rect 24 1594 26 1598
rect 30 1594 32 1598
rect 36 1594 38 1598
rect 42 1594 44 1598
rect 48 1595 64 1598
rect 68 1595 70 1599
rect 74 1595 76 1599
rect 80 1595 82 1599
rect 86 1595 89 1599
rect 93 1595 95 1599
rect 99 1595 100 1599
rect 48 1594 100 1595
rect 107 1622 135 1624
rect 111 1618 112 1622
rect 116 1618 119 1622
rect 123 1618 125 1622
rect 129 1618 131 1622
rect 107 1616 135 1618
rect 111 1612 112 1616
rect 116 1612 119 1616
rect 123 1612 125 1616
rect 129 1612 131 1616
rect 107 1610 135 1612
rect 111 1606 112 1610
rect 116 1606 119 1610
rect 123 1606 125 1610
rect 129 1606 131 1610
rect 107 1604 135 1606
rect 111 1600 112 1604
rect 116 1600 119 1604
rect 123 1600 125 1604
rect 129 1600 131 1604
rect 144 1628 148 1630
rect 144 1622 148 1624
rect 144 1616 148 1618
rect 144 1610 148 1612
rect 144 1604 148 1606
rect 107 1598 129 1600
rect 111 1594 112 1598
rect 116 1594 119 1598
rect 123 1594 125 1598
rect 144 1598 148 1600
rect 144 1592 148 1594
rect 4 1586 8 1590
rect 12 1586 63 1590
rect 72 1586 74 1590
rect 78 1586 80 1590
rect 84 1586 86 1590
rect 90 1586 92 1590
rect 101 1586 137 1590
rect 141 1588 144 1590
rect 141 1586 148 1588
rect 0 1584 144 1586
rect 4 1580 8 1584
rect 12 1580 63 1584
rect 72 1580 74 1584
rect 78 1580 80 1584
rect 84 1580 86 1584
rect 90 1580 92 1584
rect 101 1580 137 1584
rect 141 1582 144 1584
rect 141 1580 148 1582
rect 0 1578 144 1580
rect 4 1574 8 1578
rect 12 1574 63 1578
rect 72 1574 74 1578
rect 78 1574 80 1578
rect 84 1574 86 1578
rect 90 1574 92 1578
rect 101 1574 137 1578
rect 141 1576 144 1578
rect 141 1574 148 1576
rect 0 1572 144 1574
rect 4 1568 8 1572
rect 12 1568 63 1572
rect 72 1568 74 1572
rect 78 1568 80 1572
rect 84 1568 86 1572
rect 90 1568 92 1572
rect 101 1568 137 1572
rect 141 1570 144 1572
rect 141 1568 148 1570
rect 0 1566 144 1568
rect 4 1562 8 1566
rect 12 1562 63 1566
rect 72 1562 74 1566
rect 78 1562 80 1566
rect 84 1562 86 1566
rect 90 1562 92 1566
rect 101 1562 137 1566
rect 141 1564 144 1566
rect 141 1562 148 1564
rect 0 1560 144 1562
rect 4 1556 8 1560
rect 12 1556 63 1560
rect 72 1556 74 1560
rect 78 1556 80 1560
rect 84 1556 86 1560
rect 90 1556 92 1560
rect 101 1556 137 1560
rect 141 1558 144 1560
rect 141 1556 148 1558
rect 0 1554 144 1556
rect 4 1550 8 1554
rect 12 1550 63 1554
rect 72 1550 74 1554
rect 78 1550 80 1554
rect 84 1550 86 1554
rect 90 1550 92 1554
rect 101 1550 137 1554
rect 141 1552 144 1554
rect 141 1550 148 1552
rect 144 1544 148 1546
rect 144 1538 148 1540
rect 144 1532 148 1534
rect 144 1526 148 1528
rect 144 1520 148 1522
rect 144 1514 148 1516
rect 144 1508 148 1510
rect 144 1502 148 1504
rect 144 1496 148 1498
rect 144 1490 148 1492
rect 144 1484 148 1486
rect 144 1478 148 1480
rect 144 1472 148 1474
rect 144 1466 148 1468
rect 144 1460 148 1462
rect 144 1454 148 1456
rect 144 1448 148 1450
rect 144 1442 148 1444
rect 144 1436 148 1438
rect 144 1430 148 1432
rect 144 1424 148 1426
rect 148 1420 150 1424
rect 154 1420 156 1424
rect 160 1420 162 1424
rect 166 1420 168 1424
rect 172 1420 174 1424
rect 178 1420 180 1424
rect 184 1420 186 1424
rect 190 1420 192 1424
rect 196 1420 198 1424
rect 202 1420 204 1424
rect 208 1420 210 1424
rect 214 1420 216 1424
rect 220 1420 222 1424
rect 226 1420 228 1424
rect 232 1420 234 1424
rect 238 1420 240 1424
rect 244 1420 246 1424
rect 250 1420 252 1424
rect 256 1420 258 1424
rect 262 1420 264 1424
rect 268 1420 270 1424
rect 274 1420 276 1424
rect 280 1420 282 1424
rect 286 1420 288 1424
rect 292 1420 294 1424
rect 298 1420 300 1424
rect 304 1420 306 1424
rect 310 1420 312 1424
rect 316 1420 318 1424
rect 322 1420 324 1424
rect 328 1420 330 1424
rect 334 1420 336 1424
rect 340 1420 342 1424
rect 346 1420 348 1424
rect 352 1420 354 1424
rect 358 1420 360 1424
rect 364 1420 366 1424
rect 370 1420 372 1424
rect 376 1420 378 1424
rect 382 1420 384 1424
rect 388 1420 390 1424
rect 394 1420 396 1424
rect 400 1420 402 1424
rect 406 1420 408 1424
rect 412 1420 414 1424
rect 418 1420 420 1424
rect 424 1420 426 1424
rect 430 1420 432 1424
rect 436 1420 438 1424
rect 442 1420 444 1424
rect 448 1420 450 1424
rect 454 1420 456 1424
rect 460 1420 462 1424
rect 466 1420 468 1424
rect 472 1420 474 1424
rect 478 1420 480 1424
rect 484 1420 486 1424
rect 490 1420 492 1424
rect 496 1420 498 1424
rect 502 1420 504 1424
rect 508 1420 510 1424
rect 144 1418 148 1420
rect 144 1412 148 1414
rect 144 1406 148 1408
rect 144 1400 148 1402
rect 144 1394 148 1396
rect 144 1388 148 1390
rect 144 1382 148 1384
rect 144 1376 148 1378
rect 144 1370 148 1372
rect 144 1364 148 1366
rect 144 1358 148 1360
rect 144 1352 148 1354
rect 144 1346 148 1348
rect 144 1340 148 1342
rect 144 1334 148 1336
rect 144 1328 148 1330
rect 144 1322 148 1324
rect 144 1316 148 1318
rect 144 1310 148 1312
rect 144 1304 148 1306
rect 144 1298 148 1300
rect 4 1290 8 1294
rect 12 1290 63 1294
rect 72 1290 74 1294
rect 78 1290 80 1294
rect 84 1290 86 1294
rect 90 1290 92 1294
rect 101 1290 137 1294
rect 141 1292 148 1294
rect 141 1290 144 1292
rect 0 1288 144 1290
rect 4 1284 8 1288
rect 12 1284 63 1288
rect 72 1284 74 1288
rect 78 1284 80 1288
rect 84 1284 86 1288
rect 90 1284 92 1288
rect 101 1284 137 1288
rect 141 1286 148 1288
rect 141 1284 144 1286
rect 0 1282 144 1284
rect 4 1278 8 1282
rect 12 1278 63 1282
rect 72 1278 74 1282
rect 78 1278 80 1282
rect 84 1278 86 1282
rect 90 1278 92 1282
rect 101 1278 137 1282
rect 141 1280 148 1282
rect 141 1278 144 1280
rect 0 1276 144 1278
rect 4 1272 8 1276
rect 12 1272 63 1276
rect 72 1272 74 1276
rect 78 1272 80 1276
rect 84 1272 86 1276
rect 90 1272 92 1276
rect 101 1272 137 1276
rect 141 1274 148 1276
rect 141 1272 144 1274
rect 0 1270 144 1272
rect 4 1266 8 1270
rect 12 1266 63 1270
rect 72 1266 74 1270
rect 78 1266 80 1270
rect 84 1266 86 1270
rect 90 1266 92 1270
rect 101 1266 137 1270
rect 141 1268 148 1270
rect 141 1266 144 1268
rect 0 1264 144 1266
rect 4 1260 8 1264
rect 12 1260 63 1264
rect 72 1260 74 1264
rect 78 1260 80 1264
rect 84 1260 86 1264
rect 90 1260 92 1264
rect 101 1260 137 1264
rect 141 1262 148 1264
rect 141 1260 144 1262
rect 0 1258 144 1260
rect 4 1254 8 1258
rect 12 1254 63 1258
rect 72 1254 74 1258
rect 78 1254 80 1258
rect 84 1254 86 1258
rect 90 1254 92 1258
rect 101 1254 137 1258
rect 141 1256 148 1258
rect 141 1254 144 1256
rect 144 1250 148 1252
rect 4 1246 20 1250
rect 24 1246 26 1250
rect 30 1246 32 1250
rect 36 1246 38 1250
rect 42 1246 44 1250
rect 48 1249 100 1250
rect 48 1246 64 1249
rect 0 1245 64 1246
rect 68 1245 70 1249
rect 74 1245 76 1249
rect 80 1245 82 1249
rect 86 1245 89 1249
rect 93 1245 95 1249
rect 99 1245 100 1249
rect 0 1244 100 1245
rect 4 1240 14 1244
rect 18 1240 20 1244
rect 24 1240 26 1244
rect 30 1240 32 1244
rect 36 1240 38 1244
rect 42 1240 44 1244
rect 48 1243 100 1244
rect 48 1240 64 1243
rect 0 1239 64 1240
rect 68 1239 70 1243
rect 74 1239 76 1243
rect 80 1239 82 1243
rect 86 1239 89 1243
rect 93 1239 95 1243
rect 99 1239 100 1243
rect 0 1238 100 1239
rect 4 1234 14 1238
rect 18 1234 20 1238
rect 24 1234 26 1238
rect 30 1234 32 1238
rect 36 1234 38 1238
rect 42 1234 44 1238
rect 48 1237 100 1238
rect 48 1234 64 1237
rect 0 1233 64 1234
rect 68 1233 70 1237
rect 74 1233 76 1237
rect 80 1233 82 1237
rect 86 1233 89 1237
rect 93 1233 95 1237
rect 99 1233 100 1237
rect 0 1232 100 1233
rect 4 1228 14 1232
rect 18 1228 20 1232
rect 24 1228 26 1232
rect 30 1228 32 1232
rect 36 1228 38 1232
rect 42 1228 44 1232
rect 48 1231 100 1232
rect 48 1228 64 1231
rect 0 1227 64 1228
rect 68 1227 70 1231
rect 74 1227 76 1231
rect 80 1227 82 1231
rect 86 1227 89 1231
rect 93 1227 95 1231
rect 99 1227 100 1231
rect 0 1226 100 1227
rect 4 1222 14 1226
rect 18 1222 20 1226
rect 24 1222 26 1226
rect 30 1222 32 1226
rect 36 1222 38 1226
rect 42 1222 44 1226
rect 48 1225 100 1226
rect 48 1222 64 1225
rect 0 1221 64 1222
rect 68 1221 70 1225
rect 74 1221 76 1225
rect 80 1221 82 1225
rect 86 1221 89 1225
rect 93 1221 95 1225
rect 99 1221 100 1225
rect 0 1220 100 1221
rect 111 1246 112 1250
rect 116 1246 119 1250
rect 123 1246 125 1250
rect 107 1244 129 1246
rect 144 1244 148 1246
rect 111 1240 112 1244
rect 116 1240 119 1244
rect 123 1240 125 1244
rect 129 1240 131 1244
rect 107 1238 135 1240
rect 111 1234 112 1238
rect 116 1234 119 1238
rect 123 1234 125 1238
rect 129 1234 131 1238
rect 107 1232 135 1234
rect 111 1228 112 1232
rect 116 1228 119 1232
rect 123 1228 125 1232
rect 129 1228 131 1232
rect 107 1226 135 1228
rect 111 1222 112 1226
rect 116 1222 119 1226
rect 123 1222 125 1226
rect 129 1222 131 1226
rect 107 1220 135 1222
rect 4 1216 14 1220
rect 18 1216 20 1220
rect 24 1216 26 1220
rect 30 1216 32 1220
rect 36 1216 38 1220
rect 42 1216 44 1220
rect 111 1216 112 1220
rect 116 1216 119 1220
rect 123 1216 125 1220
rect 129 1216 131 1220
rect 0 1214 48 1216
rect 4 1210 14 1214
rect 18 1210 20 1214
rect 24 1210 26 1214
rect 30 1210 32 1214
rect 36 1210 38 1214
rect 42 1210 44 1214
rect 52 1212 53 1216
rect 57 1212 58 1216
rect 52 1211 58 1212
rect 52 1207 53 1211
rect 57 1207 58 1211
rect 107 1214 135 1216
rect 111 1210 112 1214
rect 116 1210 119 1214
rect 123 1210 125 1214
rect 129 1210 131 1214
rect 144 1238 148 1240
rect 144 1232 148 1234
rect 144 1226 148 1228
rect 144 1220 148 1222
rect 144 1214 148 1216
rect 52 1206 58 1207
rect 4 1202 53 1206
rect 57 1202 58 1206
rect 4 1201 58 1202
rect 4 1197 53 1201
rect 57 1197 58 1201
rect 144 1208 148 1210
rect 144 1202 148 1204
rect 4 1169 53 1173
rect 57 1169 58 1173
rect 4 1168 58 1169
rect 4 1164 53 1168
rect 57 1164 58 1168
rect 52 1163 58 1164
rect 4 1156 14 1160
rect 18 1156 20 1160
rect 24 1156 26 1160
rect 30 1156 32 1160
rect 36 1156 38 1160
rect 42 1156 44 1160
rect 0 1154 48 1156
rect 52 1159 53 1163
rect 57 1159 58 1163
rect 144 1166 148 1168
rect 144 1160 148 1162
rect 52 1158 58 1159
rect 52 1154 53 1158
rect 57 1154 58 1158
rect 111 1156 112 1160
rect 116 1156 119 1160
rect 123 1156 125 1160
rect 129 1156 131 1160
rect 107 1154 135 1156
rect 4 1150 14 1154
rect 18 1150 20 1154
rect 24 1150 26 1154
rect 30 1150 32 1154
rect 36 1150 38 1154
rect 42 1150 44 1154
rect 111 1150 112 1154
rect 116 1150 119 1154
rect 123 1150 125 1154
rect 129 1150 131 1154
rect 0 1149 100 1150
rect 0 1148 64 1149
rect 4 1144 14 1148
rect 18 1144 20 1148
rect 24 1144 26 1148
rect 30 1144 32 1148
rect 36 1144 38 1148
rect 42 1144 44 1148
rect 48 1145 64 1148
rect 68 1145 70 1149
rect 74 1145 76 1149
rect 80 1145 82 1149
rect 86 1145 89 1149
rect 93 1145 95 1149
rect 99 1145 100 1149
rect 48 1144 100 1145
rect 0 1143 100 1144
rect 0 1142 64 1143
rect 4 1138 14 1142
rect 18 1138 20 1142
rect 24 1138 26 1142
rect 30 1138 32 1142
rect 36 1138 38 1142
rect 42 1138 44 1142
rect 48 1139 64 1142
rect 68 1139 70 1143
rect 74 1139 76 1143
rect 80 1139 82 1143
rect 86 1139 89 1143
rect 93 1139 95 1143
rect 99 1139 100 1143
rect 48 1138 100 1139
rect 0 1137 100 1138
rect 0 1136 64 1137
rect 4 1132 14 1136
rect 18 1132 20 1136
rect 24 1132 26 1136
rect 30 1132 32 1136
rect 36 1132 38 1136
rect 42 1132 44 1136
rect 48 1133 64 1136
rect 68 1133 70 1137
rect 74 1133 76 1137
rect 80 1133 82 1137
rect 86 1133 89 1137
rect 93 1133 95 1137
rect 99 1133 100 1137
rect 48 1132 100 1133
rect 0 1131 100 1132
rect 0 1130 64 1131
rect 4 1126 14 1130
rect 18 1126 20 1130
rect 24 1126 26 1130
rect 30 1126 32 1130
rect 36 1126 38 1130
rect 42 1126 44 1130
rect 48 1127 64 1130
rect 68 1127 70 1131
rect 74 1127 76 1131
rect 80 1127 82 1131
rect 86 1127 89 1131
rect 93 1127 95 1131
rect 99 1127 100 1131
rect 48 1126 100 1127
rect 0 1125 100 1126
rect 0 1124 64 1125
rect 4 1120 20 1124
rect 24 1120 26 1124
rect 30 1120 32 1124
rect 36 1120 38 1124
rect 42 1120 44 1124
rect 48 1121 64 1124
rect 68 1121 70 1125
rect 74 1121 76 1125
rect 80 1121 82 1125
rect 86 1121 89 1125
rect 93 1121 95 1125
rect 99 1121 100 1125
rect 48 1120 100 1121
rect 107 1148 135 1150
rect 111 1144 112 1148
rect 116 1144 119 1148
rect 123 1144 125 1148
rect 129 1144 131 1148
rect 107 1142 135 1144
rect 111 1138 112 1142
rect 116 1138 119 1142
rect 123 1138 125 1142
rect 129 1138 131 1142
rect 107 1136 135 1138
rect 111 1132 112 1136
rect 116 1132 119 1136
rect 123 1132 125 1136
rect 129 1132 131 1136
rect 107 1130 135 1132
rect 111 1126 112 1130
rect 116 1126 119 1130
rect 123 1126 125 1130
rect 129 1126 131 1130
rect 144 1154 148 1156
rect 144 1148 148 1150
rect 144 1142 148 1144
rect 144 1136 148 1138
rect 144 1130 148 1132
rect 107 1124 129 1126
rect 111 1120 112 1124
rect 116 1120 119 1124
rect 123 1120 125 1124
rect 144 1124 148 1126
rect 144 1118 148 1120
rect 4 1112 8 1116
rect 12 1112 63 1116
rect 72 1112 74 1116
rect 78 1112 80 1116
rect 84 1112 86 1116
rect 90 1112 92 1116
rect 101 1112 137 1116
rect 141 1114 144 1116
rect 141 1112 148 1114
rect 0 1110 144 1112
rect 4 1106 8 1110
rect 12 1106 63 1110
rect 72 1106 74 1110
rect 78 1106 80 1110
rect 84 1106 86 1110
rect 90 1106 92 1110
rect 101 1106 137 1110
rect 141 1108 144 1110
rect 141 1106 148 1108
rect 0 1104 144 1106
rect 4 1100 8 1104
rect 12 1100 63 1104
rect 72 1100 74 1104
rect 78 1100 80 1104
rect 84 1100 86 1104
rect 90 1100 92 1104
rect 101 1100 137 1104
rect 141 1102 144 1104
rect 141 1100 148 1102
rect 0 1098 144 1100
rect 4 1094 8 1098
rect 12 1094 63 1098
rect 72 1094 74 1098
rect 78 1094 80 1098
rect 84 1094 86 1098
rect 90 1094 92 1098
rect 101 1094 137 1098
rect 141 1096 144 1098
rect 141 1094 148 1096
rect 0 1092 144 1094
rect 4 1088 8 1092
rect 12 1088 63 1092
rect 72 1088 74 1092
rect 78 1088 80 1092
rect 84 1088 86 1092
rect 90 1088 92 1092
rect 101 1088 137 1092
rect 141 1090 144 1092
rect 141 1088 148 1090
rect 0 1086 144 1088
rect 4 1082 8 1086
rect 12 1082 63 1086
rect 72 1082 74 1086
rect 78 1082 80 1086
rect 84 1082 86 1086
rect 90 1082 92 1086
rect 101 1082 137 1086
rect 141 1084 144 1086
rect 141 1082 148 1084
rect 0 1080 144 1082
rect 4 1076 8 1080
rect 12 1076 63 1080
rect 72 1076 74 1080
rect 78 1076 80 1080
rect 84 1076 86 1080
rect 90 1076 92 1080
rect 101 1076 137 1080
rect 141 1078 144 1080
rect 141 1076 148 1078
rect 144 1070 148 1072
rect 144 1064 148 1066
rect 144 1058 148 1060
rect 144 1052 148 1054
rect 144 1046 148 1048
rect 144 1040 148 1042
rect 144 1034 148 1036
rect 144 1028 148 1030
rect 144 1022 148 1024
rect 144 1016 148 1018
rect 144 1010 148 1012
rect 144 1004 148 1006
rect 144 998 148 1000
rect 144 992 148 994
rect 144 986 148 988
rect 144 980 148 982
rect 144 974 148 976
rect 144 968 148 970
rect 144 962 148 964
rect 144 956 148 958
rect 144 950 148 952
rect 148 946 150 950
rect 154 946 156 950
rect 160 946 162 950
rect 166 946 168 950
rect 172 946 174 950
rect 178 946 180 950
rect 184 946 186 950
rect 190 946 192 950
rect 196 946 198 950
rect 202 946 204 950
rect 208 946 210 950
rect 214 946 216 950
rect 220 946 222 950
rect 226 946 228 950
rect 232 946 234 950
rect 238 946 240 950
rect 244 946 246 950
rect 250 946 252 950
rect 256 946 258 950
rect 262 946 264 950
rect 268 946 270 950
rect 274 946 276 950
rect 280 946 282 950
rect 286 946 288 950
rect 292 946 294 950
rect 298 946 300 950
rect 304 946 306 950
rect 310 946 312 950
rect 316 946 318 950
rect 322 946 324 950
rect 328 946 330 950
rect 334 946 336 950
rect 340 946 342 950
rect 346 946 348 950
rect 352 946 354 950
rect 358 946 360 950
rect 364 946 366 950
rect 370 946 372 950
rect 376 946 378 950
rect 382 946 384 950
rect 388 946 390 950
rect 394 946 396 950
rect 400 946 402 950
rect 406 946 408 950
rect 412 946 414 950
rect 418 946 420 950
rect 424 946 426 950
rect 430 946 432 950
rect 436 946 438 950
rect 442 946 444 950
rect 448 946 450 950
rect 454 946 456 950
rect 460 946 462 950
rect 466 946 468 950
rect 472 946 474 950
rect 478 946 480 950
rect 484 946 486 950
rect 490 946 492 950
rect 496 946 498 950
rect 502 946 504 950
rect 508 946 510 950
rect 144 944 148 946
rect 144 938 148 940
rect 144 932 148 934
rect 144 926 148 928
rect 144 920 148 922
rect 144 914 148 916
rect 144 908 148 910
rect 144 902 148 904
rect 144 896 148 898
rect 144 890 148 892
rect 144 884 148 886
rect 144 878 148 880
rect 144 872 148 874
rect 144 866 148 868
rect 144 860 148 862
rect 144 854 148 856
rect 144 848 148 850
rect 144 842 148 844
rect 144 836 148 838
rect 144 830 148 832
rect 144 824 148 826
rect 4 816 8 820
rect 12 816 63 820
rect 72 816 74 820
rect 78 816 80 820
rect 84 816 86 820
rect 90 816 92 820
rect 101 816 137 820
rect 141 818 148 820
rect 141 816 144 818
rect 0 814 144 816
rect 4 810 8 814
rect 12 810 63 814
rect 72 810 74 814
rect 78 810 80 814
rect 84 810 86 814
rect 90 810 92 814
rect 101 810 137 814
rect 141 812 148 814
rect 141 810 144 812
rect 0 808 144 810
rect 4 804 8 808
rect 12 804 63 808
rect 72 804 74 808
rect 78 804 80 808
rect 84 804 86 808
rect 90 804 92 808
rect 101 804 137 808
rect 141 806 148 808
rect 141 804 144 806
rect 0 802 144 804
rect 4 798 8 802
rect 12 798 63 802
rect 72 798 74 802
rect 78 798 80 802
rect 84 798 86 802
rect 90 798 92 802
rect 101 798 137 802
rect 141 800 148 802
rect 141 798 144 800
rect 0 796 144 798
rect 4 792 8 796
rect 12 792 63 796
rect 72 792 74 796
rect 78 792 80 796
rect 84 792 86 796
rect 90 792 92 796
rect 101 792 137 796
rect 141 794 148 796
rect 141 792 144 794
rect 0 790 144 792
rect 4 786 8 790
rect 12 786 63 790
rect 72 786 74 790
rect 78 786 80 790
rect 84 786 86 790
rect 90 786 92 790
rect 101 786 137 790
rect 141 788 148 790
rect 141 786 144 788
rect 0 784 144 786
rect 4 780 8 784
rect 12 780 63 784
rect 72 780 74 784
rect 78 780 80 784
rect 84 780 86 784
rect 90 780 92 784
rect 101 780 137 784
rect 141 782 148 784
rect 141 780 144 782
rect 144 776 148 778
rect 4 772 20 776
rect 24 772 26 776
rect 30 772 32 776
rect 36 772 38 776
rect 42 772 44 776
rect 48 775 100 776
rect 48 772 64 775
rect 0 771 64 772
rect 68 771 70 775
rect 74 771 76 775
rect 80 771 82 775
rect 86 771 89 775
rect 93 771 95 775
rect 99 771 100 775
rect 0 770 100 771
rect 4 766 14 770
rect 18 766 20 770
rect 24 766 26 770
rect 30 766 32 770
rect 36 766 38 770
rect 42 766 44 770
rect 48 769 100 770
rect 48 766 64 769
rect 0 765 64 766
rect 68 765 70 769
rect 74 765 76 769
rect 80 765 82 769
rect 86 765 89 769
rect 93 765 95 769
rect 99 765 100 769
rect 0 764 100 765
rect 4 760 14 764
rect 18 760 20 764
rect 24 760 26 764
rect 30 760 32 764
rect 36 760 38 764
rect 42 760 44 764
rect 48 763 100 764
rect 48 760 64 763
rect 0 759 64 760
rect 68 759 70 763
rect 74 759 76 763
rect 80 759 82 763
rect 86 759 89 763
rect 93 759 95 763
rect 99 759 100 763
rect 0 758 100 759
rect 4 754 14 758
rect 18 754 20 758
rect 24 754 26 758
rect 30 754 32 758
rect 36 754 38 758
rect 42 754 44 758
rect 48 757 100 758
rect 48 754 64 757
rect 0 753 64 754
rect 68 753 70 757
rect 74 753 76 757
rect 80 753 82 757
rect 86 753 89 757
rect 93 753 95 757
rect 99 753 100 757
rect 0 752 100 753
rect 4 748 14 752
rect 18 748 20 752
rect 24 748 26 752
rect 30 748 32 752
rect 36 748 38 752
rect 42 748 44 752
rect 48 751 100 752
rect 48 748 64 751
rect 0 747 64 748
rect 68 747 70 751
rect 74 747 76 751
rect 80 747 82 751
rect 86 747 89 751
rect 93 747 95 751
rect 99 747 100 751
rect 0 746 100 747
rect 111 772 112 776
rect 116 772 119 776
rect 123 772 125 776
rect 107 770 129 772
rect 144 770 148 772
rect 111 766 112 770
rect 116 766 119 770
rect 123 766 125 770
rect 129 766 131 770
rect 107 764 135 766
rect 111 760 112 764
rect 116 760 119 764
rect 123 760 125 764
rect 129 760 131 764
rect 107 758 135 760
rect 111 754 112 758
rect 116 754 119 758
rect 123 754 125 758
rect 129 754 131 758
rect 107 752 135 754
rect 111 748 112 752
rect 116 748 119 752
rect 123 748 125 752
rect 129 748 131 752
rect 107 746 135 748
rect 4 742 14 746
rect 18 742 20 746
rect 24 742 26 746
rect 30 742 32 746
rect 36 742 38 746
rect 42 742 44 746
rect 111 742 112 746
rect 116 742 119 746
rect 123 742 125 746
rect 129 742 131 746
rect 0 740 48 742
rect 4 736 14 740
rect 18 736 20 740
rect 24 736 26 740
rect 30 736 32 740
rect 36 736 38 740
rect 42 736 44 740
rect 52 738 53 742
rect 57 738 58 742
rect 52 737 58 738
rect 52 733 53 737
rect 57 733 58 737
rect 107 740 135 742
rect 111 736 112 740
rect 116 736 119 740
rect 123 736 125 740
rect 129 736 131 740
rect 144 764 148 766
rect 144 758 148 760
rect 144 752 148 754
rect 144 746 148 748
rect 144 740 148 742
rect 52 732 58 733
rect 4 728 53 732
rect 57 728 58 732
rect 4 727 58 728
rect 4 723 53 727
rect 57 723 58 727
rect 144 734 148 736
rect 144 728 148 730
rect 4 695 53 699
rect 57 695 58 699
rect 4 694 58 695
rect 4 690 53 694
rect 57 690 58 694
rect 52 689 58 690
rect 4 682 14 686
rect 18 682 20 686
rect 24 682 26 686
rect 30 682 32 686
rect 36 682 38 686
rect 42 682 44 686
rect 0 680 48 682
rect 52 685 53 689
rect 57 685 58 689
rect 144 692 148 694
rect 144 686 148 688
rect 52 684 58 685
rect 52 680 53 684
rect 57 680 58 684
rect 111 682 112 686
rect 116 682 119 686
rect 123 682 125 686
rect 129 682 131 686
rect 107 680 135 682
rect 4 676 14 680
rect 18 676 20 680
rect 24 676 26 680
rect 30 676 32 680
rect 36 676 38 680
rect 42 676 44 680
rect 111 676 112 680
rect 116 676 119 680
rect 123 676 125 680
rect 129 676 131 680
rect 0 675 100 676
rect 0 674 64 675
rect 4 670 14 674
rect 18 670 20 674
rect 24 670 26 674
rect 30 670 32 674
rect 36 670 38 674
rect 42 670 44 674
rect 48 671 64 674
rect 68 671 70 675
rect 74 671 76 675
rect 80 671 82 675
rect 86 671 89 675
rect 93 671 95 675
rect 99 671 100 675
rect 48 670 100 671
rect 0 669 100 670
rect 0 668 64 669
rect 4 664 14 668
rect 18 664 20 668
rect 24 664 26 668
rect 30 664 32 668
rect 36 664 38 668
rect 42 664 44 668
rect 48 665 64 668
rect 68 665 70 669
rect 74 665 76 669
rect 80 665 82 669
rect 86 665 89 669
rect 93 665 95 669
rect 99 665 100 669
rect 48 664 100 665
rect 0 663 100 664
rect 0 662 64 663
rect 4 658 14 662
rect 18 658 20 662
rect 24 658 26 662
rect 30 658 32 662
rect 36 658 38 662
rect 42 658 44 662
rect 48 659 64 662
rect 68 659 70 663
rect 74 659 76 663
rect 80 659 82 663
rect 86 659 89 663
rect 93 659 95 663
rect 99 659 100 663
rect 48 658 100 659
rect 0 657 100 658
rect 0 656 64 657
rect 4 652 14 656
rect 18 652 20 656
rect 24 652 26 656
rect 30 652 32 656
rect 36 652 38 656
rect 42 652 44 656
rect 48 653 64 656
rect 68 653 70 657
rect 74 653 76 657
rect 80 653 82 657
rect 86 653 89 657
rect 93 653 95 657
rect 99 653 100 657
rect 48 652 100 653
rect 0 651 100 652
rect 0 650 64 651
rect 4 646 20 650
rect 24 646 26 650
rect 30 646 32 650
rect 36 646 38 650
rect 42 646 44 650
rect 48 647 64 650
rect 68 647 70 651
rect 74 647 76 651
rect 80 647 82 651
rect 86 647 89 651
rect 93 647 95 651
rect 99 647 100 651
rect 48 646 100 647
rect 107 674 135 676
rect 111 670 112 674
rect 116 670 119 674
rect 123 670 125 674
rect 129 670 131 674
rect 107 668 135 670
rect 111 664 112 668
rect 116 664 119 668
rect 123 664 125 668
rect 129 664 131 668
rect 107 662 135 664
rect 111 658 112 662
rect 116 658 119 662
rect 123 658 125 662
rect 129 658 131 662
rect 107 656 135 658
rect 111 652 112 656
rect 116 652 119 656
rect 123 652 125 656
rect 129 652 131 656
rect 144 680 148 682
rect 144 674 148 676
rect 144 668 148 670
rect 144 662 148 664
rect 144 656 148 658
rect 107 650 129 652
rect 111 646 112 650
rect 116 646 119 650
rect 123 646 125 650
rect 144 650 148 652
rect 144 644 148 646
rect 4 638 8 642
rect 12 638 63 642
rect 72 638 74 642
rect 78 638 80 642
rect 84 638 86 642
rect 90 638 92 642
rect 101 638 137 642
rect 141 640 144 642
rect 141 638 148 640
rect 0 636 144 638
rect 4 632 8 636
rect 12 632 63 636
rect 72 632 74 636
rect 78 632 80 636
rect 84 632 86 636
rect 90 632 92 636
rect 101 632 137 636
rect 141 634 144 636
rect 141 632 148 634
rect 0 630 144 632
rect 4 626 8 630
rect 12 626 63 630
rect 72 626 74 630
rect 78 626 80 630
rect 84 626 86 630
rect 90 626 92 630
rect 101 626 137 630
rect 141 628 144 630
rect 141 626 148 628
rect 0 624 144 626
rect 4 620 8 624
rect 12 620 63 624
rect 72 620 74 624
rect 78 620 80 624
rect 84 620 86 624
rect 90 620 92 624
rect 101 620 137 624
rect 141 622 144 624
rect 141 620 148 622
rect 0 618 144 620
rect 4 614 8 618
rect 12 614 63 618
rect 72 614 74 618
rect 78 614 80 618
rect 84 614 86 618
rect 90 614 92 618
rect 101 614 137 618
rect 141 616 144 618
rect 141 614 148 616
rect 0 612 144 614
rect 4 608 8 612
rect 12 608 63 612
rect 72 608 74 612
rect 78 608 80 612
rect 84 608 86 612
rect 90 608 92 612
rect 101 608 137 612
rect 141 610 144 612
rect 141 608 148 610
rect 0 606 144 608
rect 4 602 8 606
rect 12 602 63 606
rect 72 602 74 606
rect 78 602 80 606
rect 84 602 86 606
rect 90 602 92 606
rect 101 602 137 606
rect 141 604 144 606
rect 141 602 148 604
rect 144 596 148 598
rect 144 590 148 592
rect 144 584 148 586
rect 144 578 148 580
rect 144 572 148 574
rect 144 566 148 568
rect 144 560 148 562
rect 144 554 148 556
rect 144 548 148 550
rect 144 542 148 544
rect 144 536 148 538
rect 144 530 148 532
rect 144 524 148 526
rect 144 518 148 520
rect 144 512 148 514
rect 144 506 148 508
rect 144 500 148 502
rect 144 494 148 496
rect 144 488 148 490
rect 144 482 148 484
rect 144 476 148 478
rect 148 472 150 476
rect 154 472 156 476
rect 160 472 162 476
rect 166 472 168 476
rect 172 472 174 476
rect 178 472 180 476
rect 184 472 186 476
rect 190 472 192 476
rect 196 472 198 476
rect 202 472 204 476
rect 208 472 210 476
rect 214 472 216 476
rect 220 472 222 476
rect 226 472 228 476
rect 232 472 234 476
rect 238 472 240 476
rect 244 472 246 476
rect 250 472 252 476
rect 256 472 258 476
rect 262 472 264 476
rect 268 472 270 476
rect 274 472 276 476
rect 280 472 282 476
rect 286 472 288 476
rect 292 472 294 476
rect 298 472 300 476
rect 304 472 306 476
rect 310 472 312 476
rect 316 472 318 476
rect 322 472 324 476
rect 328 472 330 476
rect 334 472 336 476
rect 340 472 342 476
rect 346 472 348 476
rect 352 472 354 476
rect 358 472 360 476
rect 364 472 366 476
rect 370 472 372 476
rect 376 472 378 476
rect 382 472 384 476
rect 388 472 390 476
rect 394 472 396 476
rect 400 472 402 476
rect 406 472 408 476
rect 412 472 414 476
rect 418 472 420 476
rect 424 472 426 476
rect 430 472 432 476
rect 436 472 438 476
rect 442 472 444 476
rect 448 472 450 476
rect 454 472 456 476
rect 460 472 462 476
rect 466 472 468 476
rect 472 472 474 476
rect 478 472 480 476
rect 484 472 486 476
rect 490 472 492 476
rect 496 472 498 476
rect 502 472 504 476
rect 508 472 510 476
rect 144 470 148 472
rect 144 464 148 466
rect 144 458 148 460
rect 144 452 148 454
rect 144 446 148 448
rect 144 440 148 442
rect 144 434 148 436
rect 144 428 148 430
rect 144 422 148 424
rect 144 416 148 418
rect 144 410 148 412
rect 144 404 148 406
rect 144 398 148 400
rect 144 392 148 394
rect 144 386 148 388
rect 144 380 148 382
rect 144 374 148 376
rect 144 368 148 370
rect 144 362 148 364
rect 144 356 148 358
rect 144 350 148 352
rect 4 342 8 346
rect 12 342 63 346
rect 72 342 74 346
rect 78 342 80 346
rect 84 342 86 346
rect 90 342 92 346
rect 101 342 137 346
rect 141 344 148 346
rect 141 342 144 344
rect 0 340 144 342
rect 4 336 8 340
rect 12 336 63 340
rect 72 336 74 340
rect 78 336 80 340
rect 84 336 86 340
rect 90 336 92 340
rect 101 336 137 340
rect 141 338 148 340
rect 141 336 144 338
rect 0 334 144 336
rect 4 330 8 334
rect 12 330 63 334
rect 72 330 74 334
rect 78 330 80 334
rect 84 330 86 334
rect 90 330 92 334
rect 101 330 137 334
rect 141 332 148 334
rect 141 330 144 332
rect 0 328 144 330
rect 4 324 8 328
rect 12 324 63 328
rect 72 324 74 328
rect 78 324 80 328
rect 84 324 86 328
rect 90 324 92 328
rect 101 324 137 328
rect 141 326 148 328
rect 141 324 144 326
rect 0 322 144 324
rect 4 318 8 322
rect 12 318 63 322
rect 72 318 74 322
rect 78 318 80 322
rect 84 318 86 322
rect 90 318 92 322
rect 101 318 137 322
rect 141 320 148 322
rect 141 318 144 320
rect 0 316 144 318
rect 4 312 8 316
rect 12 312 63 316
rect 72 312 74 316
rect 78 312 80 316
rect 84 312 86 316
rect 90 312 92 316
rect 101 312 137 316
rect 141 314 148 316
rect 141 312 144 314
rect 0 310 144 312
rect 4 306 8 310
rect 12 306 63 310
rect 72 306 74 310
rect 78 306 80 310
rect 84 306 86 310
rect 90 306 92 310
rect 101 306 137 310
rect 141 308 148 310
rect 141 306 144 308
rect 144 302 148 304
rect 4 298 20 302
rect 24 298 26 302
rect 30 298 32 302
rect 36 298 38 302
rect 42 298 44 302
rect 48 301 100 302
rect 48 298 64 301
rect 0 297 64 298
rect 68 297 70 301
rect 74 297 76 301
rect 80 297 82 301
rect 86 297 89 301
rect 93 297 95 301
rect 99 297 100 301
rect 0 296 100 297
rect 4 292 14 296
rect 18 292 20 296
rect 24 292 26 296
rect 30 292 32 296
rect 36 292 38 296
rect 42 292 44 296
rect 48 295 100 296
rect 48 292 64 295
rect 0 291 64 292
rect 68 291 70 295
rect 74 291 76 295
rect 80 291 82 295
rect 86 291 89 295
rect 93 291 95 295
rect 99 291 100 295
rect 0 290 100 291
rect 4 286 14 290
rect 18 286 20 290
rect 24 286 26 290
rect 30 286 32 290
rect 36 286 38 290
rect 42 286 44 290
rect 48 289 100 290
rect 48 286 64 289
rect 0 285 64 286
rect 68 285 70 289
rect 74 285 76 289
rect 80 285 82 289
rect 86 285 89 289
rect 93 285 95 289
rect 99 285 100 289
rect 0 284 100 285
rect 4 280 14 284
rect 18 280 20 284
rect 24 280 26 284
rect 30 280 32 284
rect 36 280 38 284
rect 42 280 44 284
rect 48 283 100 284
rect 48 280 64 283
rect 0 279 64 280
rect 68 279 70 283
rect 74 279 76 283
rect 80 279 82 283
rect 86 279 89 283
rect 93 279 95 283
rect 99 279 100 283
rect 0 278 100 279
rect 4 274 14 278
rect 18 274 20 278
rect 24 274 26 278
rect 30 274 32 278
rect 36 274 38 278
rect 42 274 44 278
rect 48 277 100 278
rect 48 274 64 277
rect 0 273 64 274
rect 68 273 70 277
rect 74 273 76 277
rect 80 273 82 277
rect 86 273 89 277
rect 93 273 95 277
rect 99 273 100 277
rect 0 272 100 273
rect 111 298 112 302
rect 116 298 119 302
rect 123 298 125 302
rect 107 296 129 298
rect 144 296 148 298
rect 111 292 112 296
rect 116 292 119 296
rect 123 292 125 296
rect 129 292 131 296
rect 107 290 135 292
rect 111 286 112 290
rect 116 286 119 290
rect 123 286 125 290
rect 129 286 131 290
rect 107 284 135 286
rect 111 280 112 284
rect 116 280 119 284
rect 123 280 125 284
rect 129 280 131 284
rect 107 278 135 280
rect 111 274 112 278
rect 116 274 119 278
rect 123 274 125 278
rect 129 274 131 278
rect 107 272 135 274
rect 4 268 14 272
rect 18 268 20 272
rect 24 268 26 272
rect 30 268 32 272
rect 36 268 38 272
rect 42 268 44 272
rect 111 268 112 272
rect 116 268 119 272
rect 123 268 125 272
rect 129 268 131 272
rect 0 266 48 268
rect 4 262 14 266
rect 18 262 20 266
rect 24 262 26 266
rect 30 262 32 266
rect 36 262 38 266
rect 42 262 44 266
rect 52 264 53 268
rect 57 264 58 268
rect 52 263 58 264
rect 52 259 53 263
rect 57 259 58 263
rect 107 266 135 268
rect 111 262 112 266
rect 116 262 119 266
rect 123 262 125 266
rect 129 262 131 266
rect 144 290 148 292
rect 144 284 148 286
rect 144 278 148 280
rect 144 272 148 274
rect 144 266 148 268
rect 52 258 58 259
rect 4 254 53 258
rect 57 254 58 258
rect 4 253 58 254
rect 4 249 53 253
rect 57 249 58 253
rect 144 260 148 262
rect 144 254 148 256
rect 4 221 53 225
rect 57 221 58 225
rect 4 220 58 221
rect 4 216 53 220
rect 57 216 58 220
rect 52 215 58 216
rect 4 208 14 212
rect 18 208 20 212
rect 24 208 26 212
rect 30 208 32 212
rect 36 208 38 212
rect 42 208 44 212
rect 0 206 48 208
rect 52 211 53 215
rect 57 211 58 215
rect 144 218 148 220
rect 144 212 148 214
rect 52 210 58 211
rect 52 206 53 210
rect 57 206 58 210
rect 111 208 112 212
rect 116 208 119 212
rect 123 208 125 212
rect 129 208 131 212
rect 107 206 135 208
rect 4 202 14 206
rect 18 202 20 206
rect 24 202 26 206
rect 30 202 32 206
rect 36 202 38 206
rect 42 202 44 206
rect 111 202 112 206
rect 116 202 119 206
rect 123 202 125 206
rect 129 202 131 206
rect 0 201 100 202
rect 0 200 64 201
rect 4 196 14 200
rect 18 196 20 200
rect 24 196 26 200
rect 30 196 32 200
rect 36 196 38 200
rect 42 196 44 200
rect 48 197 64 200
rect 68 197 70 201
rect 74 197 76 201
rect 80 197 82 201
rect 86 197 89 201
rect 93 197 95 201
rect 99 197 100 201
rect 48 196 100 197
rect 0 195 100 196
rect 0 194 64 195
rect 4 190 14 194
rect 18 190 20 194
rect 24 190 26 194
rect 30 190 32 194
rect 36 190 38 194
rect 42 190 44 194
rect 48 191 64 194
rect 68 191 70 195
rect 74 191 76 195
rect 80 191 82 195
rect 86 191 89 195
rect 93 191 95 195
rect 99 191 100 195
rect 48 190 100 191
rect 0 189 100 190
rect 0 188 64 189
rect 4 184 14 188
rect 18 184 20 188
rect 24 184 26 188
rect 30 184 32 188
rect 36 184 38 188
rect 42 184 44 188
rect 48 185 64 188
rect 68 185 70 189
rect 74 185 76 189
rect 80 185 82 189
rect 86 185 89 189
rect 93 185 95 189
rect 99 185 100 189
rect 48 184 100 185
rect 0 183 100 184
rect 0 182 64 183
rect 4 178 14 182
rect 18 178 20 182
rect 24 178 26 182
rect 30 178 32 182
rect 36 178 38 182
rect 42 178 44 182
rect 48 179 64 182
rect 68 179 70 183
rect 74 179 76 183
rect 80 179 82 183
rect 86 179 89 183
rect 93 179 95 183
rect 99 179 100 183
rect 48 178 100 179
rect 0 177 100 178
rect 0 176 64 177
rect 4 172 14 176
rect 18 172 20 176
rect 24 172 26 176
rect 30 172 32 176
rect 36 172 38 176
rect 42 172 44 176
rect 48 173 64 176
rect 68 173 70 177
rect 74 173 76 177
rect 80 173 82 177
rect 86 173 89 177
rect 93 173 95 177
rect 99 173 100 177
rect 48 172 100 173
rect 107 200 135 202
rect 111 196 112 200
rect 116 196 119 200
rect 123 196 125 200
rect 129 196 131 200
rect 107 194 135 196
rect 111 190 112 194
rect 116 190 119 194
rect 123 190 125 194
rect 129 190 131 194
rect 107 188 135 190
rect 111 184 112 188
rect 116 184 119 188
rect 123 184 125 188
rect 129 184 131 188
rect 107 182 135 184
rect 111 178 112 182
rect 116 178 119 182
rect 123 178 125 182
rect 129 178 131 182
rect 144 206 148 208
rect 144 200 148 202
rect 144 194 148 196
rect 144 188 148 190
rect 144 182 148 184
rect 107 176 129 178
rect 111 172 112 176
rect 116 172 119 176
rect 123 172 125 176
rect 144 176 148 178
rect 144 170 148 172
rect 62 164 63 168
rect 72 164 74 168
rect 78 164 80 168
rect 84 164 86 168
rect 90 164 92 168
rect 101 164 137 168
rect 141 166 144 168
rect 141 164 148 166
rect 62 162 144 164
rect 62 158 63 162
rect 72 158 74 162
rect 78 158 80 162
rect 84 158 86 162
rect 90 158 92 162
rect 101 158 137 162
rect 141 160 144 162
rect 141 158 148 160
rect 62 156 144 158
rect 62 152 63 156
rect 72 152 74 156
rect 78 152 80 156
rect 84 152 86 156
rect 90 152 92 156
rect 101 152 137 156
rect 141 154 144 156
rect 141 152 148 154
rect 62 150 144 152
rect 62 146 63 150
rect 72 146 74 150
rect 78 146 80 150
rect 84 146 86 150
rect 90 146 92 150
rect 101 146 137 150
rect 141 148 144 150
rect 141 146 148 148
rect 62 144 144 146
rect 62 140 63 144
rect 72 140 74 144
rect 78 140 80 144
rect 84 140 86 144
rect 90 140 92 144
rect 101 140 137 144
rect 141 142 144 144
rect 141 140 148 142
rect 62 138 144 140
rect 62 134 63 138
rect 72 134 74 138
rect 78 134 80 138
rect 84 134 86 138
rect 90 134 92 138
rect 101 134 137 138
rect 141 136 144 138
rect 141 134 148 136
rect 62 132 144 134
rect 62 128 63 132
rect 72 128 74 132
rect 78 128 80 132
rect 84 128 86 132
rect 90 128 92 132
rect 101 128 137 132
rect 141 130 144 132
rect 141 128 148 130
rect 144 122 148 124
rect 144 116 148 118
rect 144 110 148 112
rect 144 104 148 106
rect 144 98 148 100
rect 144 92 148 94
rect 144 86 148 88
rect 144 80 148 82
rect 144 74 148 76
rect 144 68 148 70
rect 144 62 148 64
rect 144 56 148 58
rect 144 50 148 52
rect 144 44 148 46
rect 144 38 148 40
rect 144 32 148 34
rect 144 26 148 28
rect 144 20 148 22
rect 144 14 148 16
rect 144 8 148 10
rect 144 2 148 4
<< m2contact >>
rect 63 4134 72 4138
rect 74 4134 78 4138
rect 80 4134 84 4138
rect 86 4134 90 4138
rect 92 4134 101 4138
rect 63 4128 72 4132
rect 74 4128 78 4132
rect 80 4128 84 4132
rect 86 4128 90 4132
rect 92 4128 101 4132
rect 63 4122 72 4126
rect 74 4122 78 4126
rect 80 4122 84 4126
rect 86 4122 90 4126
rect 92 4122 101 4126
rect 63 4116 72 4120
rect 74 4116 78 4120
rect 80 4116 84 4120
rect 86 4116 90 4120
rect 92 4116 101 4120
rect 63 4110 72 4114
rect 74 4110 78 4114
rect 80 4110 84 4114
rect 86 4110 90 4114
rect 92 4110 101 4114
rect 63 4104 72 4108
rect 74 4104 78 4108
rect 80 4104 84 4108
rect 86 4104 90 4108
rect 92 4104 101 4108
rect 63 4098 72 4102
rect 74 4098 78 4102
rect 80 4098 84 4102
rect 86 4098 90 4102
rect 92 4098 101 4102
rect 0 4090 4 4094
rect 14 4090 18 4094
rect 26 4090 30 4094
rect 32 4090 36 4094
rect 43 4090 47 4094
rect 0 4084 4 4088
rect 14 4084 18 4088
rect 26 4084 30 4088
rect 32 4084 36 4088
rect 43 4084 47 4088
rect 0 4078 4 4082
rect 14 4078 18 4082
rect 26 4078 30 4082
rect 32 4078 36 4082
rect 43 4078 47 4082
rect 0 4072 4 4076
rect 14 4072 18 4076
rect 26 4072 30 4076
rect 32 4072 36 4076
rect 43 4072 47 4076
rect 0 4066 4 4070
rect 14 4066 18 4070
rect 26 4066 30 4070
rect 32 4066 36 4070
rect 43 4066 47 4070
rect 107 4090 111 4094
rect 119 4090 123 4094
rect 107 4084 111 4088
rect 119 4084 123 4088
rect 131 4084 135 4088
rect 107 4078 111 4082
rect 119 4078 123 4082
rect 131 4078 135 4082
rect 107 4072 111 4076
rect 119 4072 123 4076
rect 131 4072 135 4076
rect 107 4066 111 4070
rect 119 4066 123 4070
rect 131 4066 135 4070
rect 0 4060 4 4064
rect 14 4060 18 4064
rect 26 4060 30 4064
rect 32 4060 36 4064
rect 43 4060 47 4064
rect 107 4060 111 4064
rect 119 4060 123 4064
rect 131 4060 135 4064
rect 0 4054 4 4058
rect 14 4054 18 4058
rect 26 4054 30 4058
rect 32 4054 36 4058
rect 43 4054 47 4058
rect 53 4051 57 4055
rect 107 4054 111 4058
rect 119 4054 123 4058
rect 131 4054 135 4058
rect 0 4041 4 4050
rect 53 4041 57 4045
rect 0 4008 4 4017
rect 53 4013 57 4017
rect 0 4000 4 4004
rect 14 4000 18 4004
rect 26 4000 30 4004
rect 32 4000 36 4004
rect 43 4000 47 4004
rect 53 4003 57 4007
rect 107 4000 111 4004
rect 119 4000 123 4004
rect 131 4000 135 4004
rect 0 3994 4 3998
rect 14 3994 18 3998
rect 26 3994 30 3998
rect 32 3994 36 3998
rect 43 3994 47 3998
rect 107 3994 111 3998
rect 119 3994 123 3998
rect 131 3994 135 3998
rect 0 3988 4 3992
rect 14 3988 18 3992
rect 26 3988 30 3992
rect 32 3988 36 3992
rect 43 3988 47 3992
rect 0 3982 4 3986
rect 14 3982 18 3986
rect 26 3982 30 3986
rect 32 3982 36 3986
rect 43 3982 47 3986
rect 0 3976 4 3980
rect 14 3976 18 3980
rect 26 3976 30 3980
rect 32 3976 36 3980
rect 43 3976 47 3980
rect 0 3970 4 3974
rect 14 3970 18 3974
rect 26 3970 30 3974
rect 32 3970 36 3974
rect 43 3970 47 3974
rect 0 3964 4 3968
rect 26 3964 30 3968
rect 32 3964 36 3968
rect 43 3964 47 3968
rect 107 3988 111 3992
rect 119 3988 123 3992
rect 131 3988 135 3992
rect 107 3982 111 3986
rect 119 3982 123 3986
rect 131 3982 135 3986
rect 107 3976 111 3980
rect 119 3976 123 3980
rect 131 3976 135 3980
rect 107 3970 111 3974
rect 119 3970 123 3974
rect 131 3970 135 3974
rect 107 3964 111 3968
rect 119 3964 123 3968
rect 0 3956 4 3960
rect 63 3956 72 3960
rect 74 3956 78 3960
rect 80 3956 84 3960
rect 86 3956 90 3960
rect 92 3956 101 3960
rect 0 3950 4 3954
rect 63 3950 72 3954
rect 74 3950 78 3954
rect 80 3950 84 3954
rect 86 3950 90 3954
rect 92 3950 101 3954
rect 0 3944 4 3948
rect 63 3944 72 3948
rect 74 3944 78 3948
rect 80 3944 84 3948
rect 86 3944 90 3948
rect 92 3944 101 3948
rect 0 3938 4 3942
rect 63 3938 72 3942
rect 74 3938 78 3942
rect 80 3938 84 3942
rect 86 3938 90 3942
rect 92 3938 101 3942
rect 0 3932 4 3936
rect 63 3932 72 3936
rect 74 3932 78 3936
rect 80 3932 84 3936
rect 86 3932 90 3936
rect 92 3932 101 3936
rect 0 3926 4 3930
rect 63 3926 72 3930
rect 74 3926 78 3930
rect 80 3926 84 3930
rect 86 3926 90 3930
rect 92 3926 101 3930
rect 0 3920 4 3924
rect 63 3920 72 3924
rect 74 3920 78 3924
rect 80 3920 84 3924
rect 86 3920 90 3924
rect 92 3920 101 3924
rect 0 3660 4 3664
rect 63 3660 72 3664
rect 74 3660 78 3664
rect 80 3660 84 3664
rect 86 3660 90 3664
rect 92 3660 101 3664
rect 0 3654 4 3658
rect 63 3654 72 3658
rect 74 3654 78 3658
rect 80 3654 84 3658
rect 86 3654 90 3658
rect 92 3654 101 3658
rect 0 3648 4 3652
rect 63 3648 72 3652
rect 74 3648 78 3652
rect 80 3648 84 3652
rect 86 3648 90 3652
rect 92 3648 101 3652
rect 0 3642 4 3646
rect 63 3642 72 3646
rect 74 3642 78 3646
rect 80 3642 84 3646
rect 86 3642 90 3646
rect 92 3642 101 3646
rect 0 3636 4 3640
rect 63 3636 72 3640
rect 74 3636 78 3640
rect 80 3636 84 3640
rect 86 3636 90 3640
rect 92 3636 101 3640
rect 0 3630 4 3634
rect 63 3630 72 3634
rect 74 3630 78 3634
rect 80 3630 84 3634
rect 86 3630 90 3634
rect 92 3630 101 3634
rect 0 3624 4 3628
rect 63 3624 72 3628
rect 74 3624 78 3628
rect 80 3624 84 3628
rect 86 3624 90 3628
rect 92 3624 101 3628
rect 0 3616 4 3620
rect 26 3616 30 3620
rect 32 3616 36 3620
rect 44 3616 48 3620
rect 0 3610 4 3614
rect 14 3610 18 3614
rect 26 3610 30 3614
rect 32 3610 36 3614
rect 44 3610 48 3614
rect 0 3604 4 3608
rect 14 3604 18 3608
rect 26 3604 30 3608
rect 32 3604 36 3608
rect 44 3604 48 3608
rect 0 3598 4 3602
rect 14 3598 18 3602
rect 26 3598 30 3602
rect 32 3598 36 3602
rect 44 3598 48 3602
rect 0 3592 4 3596
rect 14 3592 18 3596
rect 26 3592 30 3596
rect 32 3592 36 3596
rect 44 3592 48 3596
rect 107 3616 111 3620
rect 119 3616 123 3620
rect 107 3610 111 3614
rect 119 3610 123 3614
rect 131 3610 135 3614
rect 107 3604 111 3608
rect 119 3604 123 3608
rect 131 3604 135 3608
rect 107 3598 111 3602
rect 119 3598 123 3602
rect 131 3598 135 3602
rect 107 3592 111 3596
rect 119 3592 123 3596
rect 131 3592 135 3596
rect 0 3586 4 3590
rect 14 3586 18 3590
rect 26 3586 30 3590
rect 32 3586 36 3590
rect 44 3586 48 3590
rect 107 3586 111 3590
rect 119 3586 123 3590
rect 131 3586 135 3590
rect 0 3580 4 3584
rect 14 3580 18 3584
rect 26 3580 30 3584
rect 32 3580 36 3584
rect 44 3580 48 3584
rect 53 3577 57 3581
rect 107 3580 111 3584
rect 119 3580 123 3584
rect 131 3580 135 3584
rect 0 3567 4 3576
rect 53 3567 57 3571
rect 0 3534 4 3543
rect 53 3539 57 3543
rect 0 3526 4 3530
rect 14 3526 18 3530
rect 26 3526 30 3530
rect 32 3526 36 3530
rect 44 3526 48 3530
rect 53 3529 57 3533
rect 107 3526 111 3530
rect 119 3526 123 3530
rect 131 3526 135 3530
rect 0 3520 4 3524
rect 14 3520 18 3524
rect 26 3520 30 3524
rect 32 3520 36 3524
rect 44 3520 48 3524
rect 107 3520 111 3524
rect 119 3520 123 3524
rect 131 3520 135 3524
rect 0 3514 4 3518
rect 14 3514 18 3518
rect 26 3514 30 3518
rect 32 3514 36 3518
rect 44 3514 48 3518
rect 0 3508 4 3512
rect 14 3508 18 3512
rect 26 3508 30 3512
rect 32 3508 36 3512
rect 44 3508 48 3512
rect 0 3502 4 3506
rect 14 3502 18 3506
rect 26 3502 30 3506
rect 32 3502 36 3506
rect 44 3502 48 3506
rect 0 3496 4 3500
rect 14 3496 18 3500
rect 26 3496 30 3500
rect 32 3496 36 3500
rect 44 3496 48 3500
rect 0 3490 4 3494
rect 26 3490 30 3494
rect 32 3490 36 3494
rect 44 3490 48 3494
rect 107 3514 111 3518
rect 119 3514 123 3518
rect 131 3514 135 3518
rect 107 3508 111 3512
rect 119 3508 123 3512
rect 131 3508 135 3512
rect 107 3502 111 3506
rect 119 3502 123 3506
rect 131 3502 135 3506
rect 107 3496 111 3500
rect 119 3496 123 3500
rect 131 3496 135 3500
rect 107 3490 111 3494
rect 119 3490 123 3494
rect 0 3482 4 3486
rect 63 3482 72 3486
rect 74 3482 78 3486
rect 80 3482 84 3486
rect 86 3482 90 3486
rect 92 3482 101 3486
rect 0 3476 4 3480
rect 63 3476 72 3480
rect 74 3476 78 3480
rect 80 3476 84 3480
rect 86 3476 90 3480
rect 92 3476 101 3480
rect 0 3470 4 3474
rect 63 3470 72 3474
rect 74 3470 78 3474
rect 80 3470 84 3474
rect 86 3470 90 3474
rect 92 3470 101 3474
rect 0 3464 4 3468
rect 63 3464 72 3468
rect 74 3464 78 3468
rect 80 3464 84 3468
rect 86 3464 90 3468
rect 92 3464 101 3468
rect 0 3458 4 3462
rect 63 3458 72 3462
rect 74 3458 78 3462
rect 80 3458 84 3462
rect 86 3458 90 3462
rect 92 3458 101 3462
rect 0 3452 4 3456
rect 63 3452 72 3456
rect 74 3452 78 3456
rect 80 3452 84 3456
rect 86 3452 90 3456
rect 92 3452 101 3456
rect 0 3446 4 3450
rect 63 3446 72 3450
rect 74 3446 78 3450
rect 80 3446 84 3450
rect 86 3446 90 3450
rect 92 3446 101 3450
rect 0 3186 4 3190
rect 63 3186 72 3190
rect 74 3186 78 3190
rect 80 3186 84 3190
rect 86 3186 90 3190
rect 92 3186 101 3190
rect 0 3180 4 3184
rect 63 3180 72 3184
rect 74 3180 78 3184
rect 80 3180 84 3184
rect 86 3180 90 3184
rect 92 3180 101 3184
rect 0 3174 4 3178
rect 63 3174 72 3178
rect 74 3174 78 3178
rect 80 3174 84 3178
rect 86 3174 90 3178
rect 92 3174 101 3178
rect 0 3168 4 3172
rect 63 3168 72 3172
rect 74 3168 78 3172
rect 80 3168 84 3172
rect 86 3168 90 3172
rect 92 3168 101 3172
rect 0 3162 4 3166
rect 63 3162 72 3166
rect 74 3162 78 3166
rect 80 3162 84 3166
rect 86 3162 90 3166
rect 92 3162 101 3166
rect 0 3156 4 3160
rect 63 3156 72 3160
rect 74 3156 78 3160
rect 80 3156 84 3160
rect 86 3156 90 3160
rect 92 3156 101 3160
rect 0 3150 4 3154
rect 63 3150 72 3154
rect 74 3150 78 3154
rect 80 3150 84 3154
rect 86 3150 90 3154
rect 92 3150 101 3154
rect 0 3142 4 3146
rect 26 3142 30 3146
rect 32 3142 36 3146
rect 44 3142 48 3146
rect 0 3136 4 3140
rect 14 3136 18 3140
rect 26 3136 30 3140
rect 32 3136 36 3140
rect 44 3136 48 3140
rect 0 3130 4 3134
rect 14 3130 18 3134
rect 26 3130 30 3134
rect 32 3130 36 3134
rect 44 3130 48 3134
rect 0 3124 4 3128
rect 14 3124 18 3128
rect 26 3124 30 3128
rect 32 3124 36 3128
rect 44 3124 48 3128
rect 0 3118 4 3122
rect 14 3118 18 3122
rect 26 3118 30 3122
rect 32 3118 36 3122
rect 44 3118 48 3122
rect 107 3142 111 3146
rect 119 3142 123 3146
rect 107 3136 111 3140
rect 119 3136 123 3140
rect 131 3136 135 3140
rect 107 3130 111 3134
rect 119 3130 123 3134
rect 131 3130 135 3134
rect 107 3124 111 3128
rect 119 3124 123 3128
rect 131 3124 135 3128
rect 107 3118 111 3122
rect 119 3118 123 3122
rect 131 3118 135 3122
rect 0 3112 4 3116
rect 14 3112 18 3116
rect 26 3112 30 3116
rect 32 3112 36 3116
rect 44 3112 48 3116
rect 107 3112 111 3116
rect 119 3112 123 3116
rect 131 3112 135 3116
rect 0 3106 4 3110
rect 14 3106 18 3110
rect 26 3106 30 3110
rect 32 3106 36 3110
rect 44 3106 48 3110
rect 53 3103 57 3107
rect 107 3106 111 3110
rect 119 3106 123 3110
rect 131 3106 135 3110
rect 0 3093 4 3102
rect 53 3093 57 3097
rect 0 3060 4 3069
rect 53 3065 57 3069
rect 0 3052 4 3056
rect 14 3052 18 3056
rect 26 3052 30 3056
rect 32 3052 36 3056
rect 44 3052 48 3056
rect 53 3055 57 3059
rect 107 3052 111 3056
rect 119 3052 123 3056
rect 131 3052 135 3056
rect 0 3046 4 3050
rect 14 3046 18 3050
rect 26 3046 30 3050
rect 32 3046 36 3050
rect 44 3046 48 3050
rect 107 3046 111 3050
rect 119 3046 123 3050
rect 131 3046 135 3050
rect 0 3040 4 3044
rect 14 3040 18 3044
rect 26 3040 30 3044
rect 32 3040 36 3044
rect 44 3040 48 3044
rect 0 3034 4 3038
rect 14 3034 18 3038
rect 26 3034 30 3038
rect 32 3034 36 3038
rect 44 3034 48 3038
rect 0 3028 4 3032
rect 14 3028 18 3032
rect 26 3028 30 3032
rect 32 3028 36 3032
rect 44 3028 48 3032
rect 0 3022 4 3026
rect 14 3022 18 3026
rect 26 3022 30 3026
rect 32 3022 36 3026
rect 44 3022 48 3026
rect 0 3016 4 3020
rect 26 3016 30 3020
rect 32 3016 36 3020
rect 44 3016 48 3020
rect 107 3040 111 3044
rect 119 3040 123 3044
rect 131 3040 135 3044
rect 107 3034 111 3038
rect 119 3034 123 3038
rect 131 3034 135 3038
rect 107 3028 111 3032
rect 119 3028 123 3032
rect 131 3028 135 3032
rect 107 3022 111 3026
rect 119 3022 123 3026
rect 131 3022 135 3026
rect 107 3016 111 3020
rect 119 3016 123 3020
rect 0 3008 4 3012
rect 63 3008 72 3012
rect 74 3008 78 3012
rect 80 3008 84 3012
rect 86 3008 90 3012
rect 92 3008 101 3012
rect 0 3002 4 3006
rect 63 3002 72 3006
rect 74 3002 78 3006
rect 80 3002 84 3006
rect 86 3002 90 3006
rect 92 3002 101 3006
rect 0 2996 4 3000
rect 63 2996 72 3000
rect 74 2996 78 3000
rect 80 2996 84 3000
rect 86 2996 90 3000
rect 92 2996 101 3000
rect 0 2990 4 2994
rect 63 2990 72 2994
rect 74 2990 78 2994
rect 80 2990 84 2994
rect 86 2990 90 2994
rect 92 2990 101 2994
rect 0 2984 4 2988
rect 63 2984 72 2988
rect 74 2984 78 2988
rect 80 2984 84 2988
rect 86 2984 90 2988
rect 92 2984 101 2988
rect 0 2978 4 2982
rect 63 2978 72 2982
rect 74 2978 78 2982
rect 80 2978 84 2982
rect 86 2978 90 2982
rect 92 2978 101 2982
rect 0 2972 4 2976
rect 63 2972 72 2976
rect 74 2972 78 2976
rect 80 2972 84 2976
rect 86 2972 90 2976
rect 92 2972 101 2976
rect 0 2712 4 2716
rect 63 2712 72 2716
rect 74 2712 78 2716
rect 80 2712 84 2716
rect 86 2712 90 2716
rect 92 2712 101 2716
rect 0 2706 4 2710
rect 63 2706 72 2710
rect 74 2706 78 2710
rect 80 2706 84 2710
rect 86 2706 90 2710
rect 92 2706 101 2710
rect 0 2700 4 2704
rect 63 2700 72 2704
rect 74 2700 78 2704
rect 80 2700 84 2704
rect 86 2700 90 2704
rect 92 2700 101 2704
rect 0 2694 4 2698
rect 63 2694 72 2698
rect 74 2694 78 2698
rect 80 2694 84 2698
rect 86 2694 90 2698
rect 92 2694 101 2698
rect 0 2688 4 2692
rect 63 2688 72 2692
rect 74 2688 78 2692
rect 80 2688 84 2692
rect 86 2688 90 2692
rect 92 2688 101 2692
rect 0 2682 4 2686
rect 63 2682 72 2686
rect 74 2682 78 2686
rect 80 2682 84 2686
rect 86 2682 90 2686
rect 92 2682 101 2686
rect 0 2676 4 2680
rect 63 2676 72 2680
rect 74 2676 78 2680
rect 80 2676 84 2680
rect 86 2676 90 2680
rect 92 2676 101 2680
rect 0 2668 4 2672
rect 26 2668 30 2672
rect 32 2668 36 2672
rect 44 2668 48 2672
rect 0 2662 4 2666
rect 14 2662 18 2666
rect 26 2662 30 2666
rect 32 2662 36 2666
rect 44 2662 48 2666
rect 0 2656 4 2660
rect 14 2656 18 2660
rect 26 2656 30 2660
rect 32 2656 36 2660
rect 44 2656 48 2660
rect 0 2650 4 2654
rect 14 2650 18 2654
rect 26 2650 30 2654
rect 32 2650 36 2654
rect 44 2650 48 2654
rect 0 2644 4 2648
rect 14 2644 18 2648
rect 26 2644 30 2648
rect 32 2644 36 2648
rect 44 2644 48 2648
rect 107 2668 111 2672
rect 119 2668 123 2672
rect 107 2662 111 2666
rect 119 2662 123 2666
rect 131 2662 135 2666
rect 107 2656 111 2660
rect 119 2656 123 2660
rect 131 2656 135 2660
rect 107 2650 111 2654
rect 119 2650 123 2654
rect 131 2650 135 2654
rect 107 2644 111 2648
rect 119 2644 123 2648
rect 131 2644 135 2648
rect 0 2638 4 2642
rect 14 2638 18 2642
rect 26 2638 30 2642
rect 32 2638 36 2642
rect 44 2638 48 2642
rect 107 2638 111 2642
rect 119 2638 123 2642
rect 131 2638 135 2642
rect 0 2632 4 2636
rect 14 2632 18 2636
rect 26 2632 30 2636
rect 32 2632 36 2636
rect 44 2632 48 2636
rect 53 2629 57 2633
rect 107 2632 111 2636
rect 119 2632 123 2636
rect 131 2632 135 2636
rect 0 2619 4 2628
rect 53 2619 57 2623
rect 0 2586 4 2595
rect 53 2591 57 2595
rect 0 2578 4 2582
rect 14 2578 18 2582
rect 26 2578 30 2582
rect 32 2578 36 2582
rect 44 2578 48 2582
rect 53 2581 57 2585
rect 107 2578 111 2582
rect 119 2578 123 2582
rect 131 2578 135 2582
rect 0 2572 4 2576
rect 14 2572 18 2576
rect 26 2572 30 2576
rect 32 2572 36 2576
rect 44 2572 48 2576
rect 107 2572 111 2576
rect 119 2572 123 2576
rect 131 2572 135 2576
rect 0 2566 4 2570
rect 14 2566 18 2570
rect 26 2566 30 2570
rect 32 2566 36 2570
rect 44 2566 48 2570
rect 0 2560 4 2564
rect 14 2560 18 2564
rect 26 2560 30 2564
rect 32 2560 36 2564
rect 44 2560 48 2564
rect 0 2554 4 2558
rect 14 2554 18 2558
rect 26 2554 30 2558
rect 32 2554 36 2558
rect 44 2554 48 2558
rect 0 2548 4 2552
rect 14 2548 18 2552
rect 26 2548 30 2552
rect 32 2548 36 2552
rect 44 2548 48 2552
rect 0 2542 4 2546
rect 26 2542 30 2546
rect 32 2542 36 2546
rect 44 2542 48 2546
rect 107 2566 111 2570
rect 119 2566 123 2570
rect 131 2566 135 2570
rect 107 2560 111 2564
rect 119 2560 123 2564
rect 131 2560 135 2564
rect 107 2554 111 2558
rect 119 2554 123 2558
rect 131 2554 135 2558
rect 107 2548 111 2552
rect 119 2548 123 2552
rect 131 2548 135 2552
rect 107 2542 111 2546
rect 119 2542 123 2546
rect 0 2534 4 2538
rect 63 2534 72 2538
rect 74 2534 78 2538
rect 80 2534 84 2538
rect 86 2534 90 2538
rect 92 2534 101 2538
rect 0 2528 4 2532
rect 63 2528 72 2532
rect 74 2528 78 2532
rect 80 2528 84 2532
rect 86 2528 90 2532
rect 92 2528 101 2532
rect 0 2522 4 2526
rect 63 2522 72 2526
rect 74 2522 78 2526
rect 80 2522 84 2526
rect 86 2522 90 2526
rect 92 2522 101 2526
rect 0 2516 4 2520
rect 63 2516 72 2520
rect 74 2516 78 2520
rect 80 2516 84 2520
rect 86 2516 90 2520
rect 92 2516 101 2520
rect 0 2510 4 2514
rect 63 2510 72 2514
rect 74 2510 78 2514
rect 80 2510 84 2514
rect 86 2510 90 2514
rect 92 2510 101 2514
rect 0 2504 4 2508
rect 63 2504 72 2508
rect 74 2504 78 2508
rect 80 2504 84 2508
rect 86 2504 90 2508
rect 92 2504 101 2508
rect 0 2498 4 2502
rect 63 2498 72 2502
rect 74 2498 78 2502
rect 80 2498 84 2502
rect 86 2498 90 2502
rect 92 2498 101 2502
rect 0 2238 4 2242
rect 63 2238 72 2242
rect 74 2238 78 2242
rect 80 2238 84 2242
rect 86 2238 90 2242
rect 92 2238 101 2242
rect 0 2232 4 2236
rect 63 2232 72 2236
rect 74 2232 78 2236
rect 80 2232 84 2236
rect 86 2232 90 2236
rect 92 2232 101 2236
rect 0 2226 4 2230
rect 63 2226 72 2230
rect 74 2226 78 2230
rect 80 2226 84 2230
rect 86 2226 90 2230
rect 92 2226 101 2230
rect 0 2220 4 2224
rect 63 2220 72 2224
rect 74 2220 78 2224
rect 80 2220 84 2224
rect 86 2220 90 2224
rect 92 2220 101 2224
rect 0 2214 4 2218
rect 63 2214 72 2218
rect 74 2214 78 2218
rect 80 2214 84 2218
rect 86 2214 90 2218
rect 92 2214 101 2218
rect 0 2208 4 2212
rect 63 2208 72 2212
rect 74 2208 78 2212
rect 80 2208 84 2212
rect 86 2208 90 2212
rect 92 2208 101 2212
rect 0 2202 4 2206
rect 63 2202 72 2206
rect 74 2202 78 2206
rect 80 2202 84 2206
rect 86 2202 90 2206
rect 92 2202 101 2206
rect 0 2194 4 2198
rect 26 2194 30 2198
rect 32 2194 36 2198
rect 44 2194 48 2198
rect 0 2188 4 2192
rect 14 2188 18 2192
rect 26 2188 30 2192
rect 32 2188 36 2192
rect 44 2188 48 2192
rect 0 2182 4 2186
rect 14 2182 18 2186
rect 26 2182 30 2186
rect 32 2182 36 2186
rect 44 2182 48 2186
rect 0 2176 4 2180
rect 14 2176 18 2180
rect 26 2176 30 2180
rect 32 2176 36 2180
rect 44 2176 48 2180
rect 0 2170 4 2174
rect 14 2170 18 2174
rect 26 2170 30 2174
rect 32 2170 36 2174
rect 44 2170 48 2174
rect 107 2194 111 2198
rect 119 2194 123 2198
rect 107 2188 111 2192
rect 119 2188 123 2192
rect 131 2188 135 2192
rect 107 2182 111 2186
rect 119 2182 123 2186
rect 131 2182 135 2186
rect 107 2176 111 2180
rect 119 2176 123 2180
rect 131 2176 135 2180
rect 107 2170 111 2174
rect 119 2170 123 2174
rect 131 2170 135 2174
rect 0 2164 4 2168
rect 14 2164 18 2168
rect 26 2164 30 2168
rect 32 2164 36 2168
rect 44 2164 48 2168
rect 107 2164 111 2168
rect 119 2164 123 2168
rect 131 2164 135 2168
rect 0 2158 4 2162
rect 14 2158 18 2162
rect 26 2158 30 2162
rect 32 2158 36 2162
rect 44 2158 48 2162
rect 53 2155 57 2159
rect 107 2158 111 2162
rect 119 2158 123 2162
rect 131 2158 135 2162
rect 0 2145 4 2154
rect 53 2145 57 2149
rect 0 2112 4 2121
rect 53 2117 57 2121
rect 0 2104 4 2108
rect 14 2104 18 2108
rect 26 2104 30 2108
rect 32 2104 36 2108
rect 44 2104 48 2108
rect 53 2107 57 2111
rect 107 2104 111 2108
rect 119 2104 123 2108
rect 131 2104 135 2108
rect 0 2098 4 2102
rect 14 2098 18 2102
rect 26 2098 30 2102
rect 32 2098 36 2102
rect 44 2098 48 2102
rect 107 2098 111 2102
rect 119 2098 123 2102
rect 131 2098 135 2102
rect 0 2092 4 2096
rect 14 2092 18 2096
rect 26 2092 30 2096
rect 32 2092 36 2096
rect 44 2092 48 2096
rect 0 2086 4 2090
rect 14 2086 18 2090
rect 26 2086 30 2090
rect 32 2086 36 2090
rect 44 2086 48 2090
rect 0 2080 4 2084
rect 14 2080 18 2084
rect 26 2080 30 2084
rect 32 2080 36 2084
rect 44 2080 48 2084
rect 0 2074 4 2078
rect 14 2074 18 2078
rect 26 2074 30 2078
rect 32 2074 36 2078
rect 44 2074 48 2078
rect 0 2068 4 2072
rect 26 2068 30 2072
rect 32 2068 36 2072
rect 44 2068 48 2072
rect 107 2092 111 2096
rect 119 2092 123 2096
rect 131 2092 135 2096
rect 107 2086 111 2090
rect 119 2086 123 2090
rect 131 2086 135 2090
rect 107 2080 111 2084
rect 119 2080 123 2084
rect 131 2080 135 2084
rect 107 2074 111 2078
rect 119 2074 123 2078
rect 131 2074 135 2078
rect 107 2068 111 2072
rect 119 2068 123 2072
rect 0 2060 4 2064
rect 63 2060 72 2064
rect 74 2060 78 2064
rect 80 2060 84 2064
rect 86 2060 90 2064
rect 92 2060 101 2064
rect 0 2054 4 2058
rect 63 2054 72 2058
rect 74 2054 78 2058
rect 80 2054 84 2058
rect 86 2054 90 2058
rect 92 2054 101 2058
rect 0 2048 4 2052
rect 63 2048 72 2052
rect 74 2048 78 2052
rect 80 2048 84 2052
rect 86 2048 90 2052
rect 92 2048 101 2052
rect 0 2042 4 2046
rect 63 2042 72 2046
rect 74 2042 78 2046
rect 80 2042 84 2046
rect 86 2042 90 2046
rect 92 2042 101 2046
rect 0 2036 4 2040
rect 63 2036 72 2040
rect 74 2036 78 2040
rect 80 2036 84 2040
rect 86 2036 90 2040
rect 92 2036 101 2040
rect 0 2030 4 2034
rect 63 2030 72 2034
rect 74 2030 78 2034
rect 80 2030 84 2034
rect 86 2030 90 2034
rect 92 2030 101 2034
rect 0 2024 4 2028
rect 63 2024 72 2028
rect 74 2024 78 2028
rect 80 2024 84 2028
rect 86 2024 90 2028
rect 92 2024 101 2028
rect 0 1764 4 1768
rect 63 1764 72 1768
rect 74 1764 78 1768
rect 80 1764 84 1768
rect 86 1764 90 1768
rect 92 1764 101 1768
rect 0 1758 4 1762
rect 63 1758 72 1762
rect 74 1758 78 1762
rect 80 1758 84 1762
rect 86 1758 90 1762
rect 92 1758 101 1762
rect 0 1752 4 1756
rect 63 1752 72 1756
rect 74 1752 78 1756
rect 80 1752 84 1756
rect 86 1752 90 1756
rect 92 1752 101 1756
rect 0 1746 4 1750
rect 63 1746 72 1750
rect 74 1746 78 1750
rect 80 1746 84 1750
rect 86 1746 90 1750
rect 92 1746 101 1750
rect 0 1740 4 1744
rect 63 1740 72 1744
rect 74 1740 78 1744
rect 80 1740 84 1744
rect 86 1740 90 1744
rect 92 1740 101 1744
rect 0 1734 4 1738
rect 63 1734 72 1738
rect 74 1734 78 1738
rect 80 1734 84 1738
rect 86 1734 90 1738
rect 92 1734 101 1738
rect 0 1728 4 1732
rect 63 1728 72 1732
rect 74 1728 78 1732
rect 80 1728 84 1732
rect 86 1728 90 1732
rect 92 1728 101 1732
rect 0 1720 4 1724
rect 26 1720 30 1724
rect 32 1720 36 1724
rect 44 1720 48 1724
rect 0 1714 4 1718
rect 14 1714 18 1718
rect 26 1714 30 1718
rect 32 1714 36 1718
rect 44 1714 48 1718
rect 0 1708 4 1712
rect 14 1708 18 1712
rect 26 1708 30 1712
rect 32 1708 36 1712
rect 44 1708 48 1712
rect 0 1702 4 1706
rect 14 1702 18 1706
rect 26 1702 30 1706
rect 32 1702 36 1706
rect 44 1702 48 1706
rect 0 1696 4 1700
rect 14 1696 18 1700
rect 26 1696 30 1700
rect 32 1696 36 1700
rect 44 1696 48 1700
rect 107 1720 111 1724
rect 119 1720 123 1724
rect 107 1714 111 1718
rect 119 1714 123 1718
rect 131 1714 135 1718
rect 107 1708 111 1712
rect 119 1708 123 1712
rect 131 1708 135 1712
rect 107 1702 111 1706
rect 119 1702 123 1706
rect 131 1702 135 1706
rect 107 1696 111 1700
rect 119 1696 123 1700
rect 131 1696 135 1700
rect 0 1690 4 1694
rect 14 1690 18 1694
rect 26 1690 30 1694
rect 32 1690 36 1694
rect 44 1690 48 1694
rect 107 1690 111 1694
rect 119 1690 123 1694
rect 131 1690 135 1694
rect 0 1684 4 1688
rect 14 1684 18 1688
rect 26 1684 30 1688
rect 32 1684 36 1688
rect 44 1684 48 1688
rect 53 1681 57 1685
rect 107 1684 111 1688
rect 119 1684 123 1688
rect 131 1684 135 1688
rect 0 1671 4 1680
rect 53 1671 57 1675
rect 0 1638 4 1647
rect 53 1643 57 1647
rect 0 1630 4 1634
rect 14 1630 18 1634
rect 26 1630 30 1634
rect 32 1630 36 1634
rect 44 1630 48 1634
rect 53 1633 57 1637
rect 107 1630 111 1634
rect 119 1630 123 1634
rect 131 1630 135 1634
rect 0 1624 4 1628
rect 14 1624 18 1628
rect 26 1624 30 1628
rect 32 1624 36 1628
rect 44 1624 48 1628
rect 107 1624 111 1628
rect 119 1624 123 1628
rect 131 1624 135 1628
rect 0 1618 4 1622
rect 14 1618 18 1622
rect 26 1618 30 1622
rect 32 1618 36 1622
rect 44 1618 48 1622
rect 0 1612 4 1616
rect 14 1612 18 1616
rect 26 1612 30 1616
rect 32 1612 36 1616
rect 44 1612 48 1616
rect 0 1606 4 1610
rect 14 1606 18 1610
rect 26 1606 30 1610
rect 32 1606 36 1610
rect 44 1606 48 1610
rect 0 1600 4 1604
rect 14 1600 18 1604
rect 26 1600 30 1604
rect 32 1600 36 1604
rect 44 1600 48 1604
rect 0 1594 4 1598
rect 26 1594 30 1598
rect 32 1594 36 1598
rect 44 1594 48 1598
rect 107 1618 111 1622
rect 119 1618 123 1622
rect 131 1618 135 1622
rect 107 1612 111 1616
rect 119 1612 123 1616
rect 131 1612 135 1616
rect 107 1606 111 1610
rect 119 1606 123 1610
rect 131 1606 135 1610
rect 107 1600 111 1604
rect 119 1600 123 1604
rect 131 1600 135 1604
rect 107 1594 111 1598
rect 119 1594 123 1598
rect 0 1586 4 1590
rect 63 1586 72 1590
rect 74 1586 78 1590
rect 80 1586 84 1590
rect 86 1586 90 1590
rect 92 1586 101 1590
rect 0 1580 4 1584
rect 63 1580 72 1584
rect 74 1580 78 1584
rect 80 1580 84 1584
rect 86 1580 90 1584
rect 92 1580 101 1584
rect 0 1574 4 1578
rect 63 1574 72 1578
rect 74 1574 78 1578
rect 80 1574 84 1578
rect 86 1574 90 1578
rect 92 1574 101 1578
rect 0 1568 4 1572
rect 63 1568 72 1572
rect 74 1568 78 1572
rect 80 1568 84 1572
rect 86 1568 90 1572
rect 92 1568 101 1572
rect 0 1562 4 1566
rect 63 1562 72 1566
rect 74 1562 78 1566
rect 80 1562 84 1566
rect 86 1562 90 1566
rect 92 1562 101 1566
rect 0 1556 4 1560
rect 63 1556 72 1560
rect 74 1556 78 1560
rect 80 1556 84 1560
rect 86 1556 90 1560
rect 92 1556 101 1560
rect 0 1550 4 1554
rect 63 1550 72 1554
rect 74 1550 78 1554
rect 80 1550 84 1554
rect 86 1550 90 1554
rect 92 1550 101 1554
rect 0 1290 4 1294
rect 63 1290 72 1294
rect 74 1290 78 1294
rect 80 1290 84 1294
rect 86 1290 90 1294
rect 92 1290 101 1294
rect 0 1284 4 1288
rect 63 1284 72 1288
rect 74 1284 78 1288
rect 80 1284 84 1288
rect 86 1284 90 1288
rect 92 1284 101 1288
rect 0 1278 4 1282
rect 63 1278 72 1282
rect 74 1278 78 1282
rect 80 1278 84 1282
rect 86 1278 90 1282
rect 92 1278 101 1282
rect 0 1272 4 1276
rect 63 1272 72 1276
rect 74 1272 78 1276
rect 80 1272 84 1276
rect 86 1272 90 1276
rect 92 1272 101 1276
rect 0 1266 4 1270
rect 63 1266 72 1270
rect 74 1266 78 1270
rect 80 1266 84 1270
rect 86 1266 90 1270
rect 92 1266 101 1270
rect 0 1260 4 1264
rect 63 1260 72 1264
rect 74 1260 78 1264
rect 80 1260 84 1264
rect 86 1260 90 1264
rect 92 1260 101 1264
rect 0 1254 4 1258
rect 63 1254 72 1258
rect 74 1254 78 1258
rect 80 1254 84 1258
rect 86 1254 90 1258
rect 92 1254 101 1258
rect 0 1246 4 1250
rect 26 1246 30 1250
rect 32 1246 36 1250
rect 44 1246 48 1250
rect 0 1240 4 1244
rect 14 1240 18 1244
rect 26 1240 30 1244
rect 32 1240 36 1244
rect 44 1240 48 1244
rect 0 1234 4 1238
rect 14 1234 18 1238
rect 26 1234 30 1238
rect 32 1234 36 1238
rect 44 1234 48 1238
rect 0 1228 4 1232
rect 14 1228 18 1232
rect 26 1228 30 1232
rect 32 1228 36 1232
rect 44 1228 48 1232
rect 0 1222 4 1226
rect 14 1222 18 1226
rect 26 1222 30 1226
rect 32 1222 36 1226
rect 44 1222 48 1226
rect 107 1246 111 1250
rect 119 1246 123 1250
rect 107 1240 111 1244
rect 119 1240 123 1244
rect 131 1240 135 1244
rect 107 1234 111 1238
rect 119 1234 123 1238
rect 131 1234 135 1238
rect 107 1228 111 1232
rect 119 1228 123 1232
rect 131 1228 135 1232
rect 107 1222 111 1226
rect 119 1222 123 1226
rect 131 1222 135 1226
rect 0 1216 4 1220
rect 14 1216 18 1220
rect 26 1216 30 1220
rect 32 1216 36 1220
rect 44 1216 48 1220
rect 107 1216 111 1220
rect 119 1216 123 1220
rect 131 1216 135 1220
rect 0 1210 4 1214
rect 14 1210 18 1214
rect 26 1210 30 1214
rect 32 1210 36 1214
rect 44 1210 48 1214
rect 53 1207 57 1211
rect 107 1210 111 1214
rect 119 1210 123 1214
rect 131 1210 135 1214
rect 0 1197 4 1206
rect 53 1197 57 1201
rect 0 1164 4 1173
rect 53 1169 57 1173
rect 0 1156 4 1160
rect 14 1156 18 1160
rect 26 1156 30 1160
rect 32 1156 36 1160
rect 44 1156 48 1160
rect 53 1159 57 1163
rect 107 1156 111 1160
rect 119 1156 123 1160
rect 131 1156 135 1160
rect 0 1150 4 1154
rect 14 1150 18 1154
rect 26 1150 30 1154
rect 32 1150 36 1154
rect 44 1150 48 1154
rect 107 1150 111 1154
rect 119 1150 123 1154
rect 131 1150 135 1154
rect 0 1144 4 1148
rect 14 1144 18 1148
rect 26 1144 30 1148
rect 32 1144 36 1148
rect 44 1144 48 1148
rect 0 1138 4 1142
rect 14 1138 18 1142
rect 26 1138 30 1142
rect 32 1138 36 1142
rect 44 1138 48 1142
rect 0 1132 4 1136
rect 14 1132 18 1136
rect 26 1132 30 1136
rect 32 1132 36 1136
rect 44 1132 48 1136
rect 0 1126 4 1130
rect 14 1126 18 1130
rect 26 1126 30 1130
rect 32 1126 36 1130
rect 44 1126 48 1130
rect 0 1120 4 1124
rect 26 1120 30 1124
rect 32 1120 36 1124
rect 44 1120 48 1124
rect 107 1144 111 1148
rect 119 1144 123 1148
rect 131 1144 135 1148
rect 107 1138 111 1142
rect 119 1138 123 1142
rect 131 1138 135 1142
rect 107 1132 111 1136
rect 119 1132 123 1136
rect 131 1132 135 1136
rect 107 1126 111 1130
rect 119 1126 123 1130
rect 131 1126 135 1130
rect 107 1120 111 1124
rect 119 1120 123 1124
rect 0 1112 4 1116
rect 63 1112 72 1116
rect 74 1112 78 1116
rect 80 1112 84 1116
rect 86 1112 90 1116
rect 92 1112 101 1116
rect 0 1106 4 1110
rect 63 1106 72 1110
rect 74 1106 78 1110
rect 80 1106 84 1110
rect 86 1106 90 1110
rect 92 1106 101 1110
rect 0 1100 4 1104
rect 63 1100 72 1104
rect 74 1100 78 1104
rect 80 1100 84 1104
rect 86 1100 90 1104
rect 92 1100 101 1104
rect 0 1094 4 1098
rect 63 1094 72 1098
rect 74 1094 78 1098
rect 80 1094 84 1098
rect 86 1094 90 1098
rect 92 1094 101 1098
rect 0 1088 4 1092
rect 63 1088 72 1092
rect 74 1088 78 1092
rect 80 1088 84 1092
rect 86 1088 90 1092
rect 92 1088 101 1092
rect 0 1082 4 1086
rect 63 1082 72 1086
rect 74 1082 78 1086
rect 80 1082 84 1086
rect 86 1082 90 1086
rect 92 1082 101 1086
rect 0 1076 4 1080
rect 63 1076 72 1080
rect 74 1076 78 1080
rect 80 1076 84 1080
rect 86 1076 90 1080
rect 92 1076 101 1080
rect 0 816 4 820
rect 63 816 72 820
rect 74 816 78 820
rect 80 816 84 820
rect 86 816 90 820
rect 92 816 101 820
rect 0 810 4 814
rect 63 810 72 814
rect 74 810 78 814
rect 80 810 84 814
rect 86 810 90 814
rect 92 810 101 814
rect 0 804 4 808
rect 63 804 72 808
rect 74 804 78 808
rect 80 804 84 808
rect 86 804 90 808
rect 92 804 101 808
rect 0 798 4 802
rect 63 798 72 802
rect 74 798 78 802
rect 80 798 84 802
rect 86 798 90 802
rect 92 798 101 802
rect 0 792 4 796
rect 63 792 72 796
rect 74 792 78 796
rect 80 792 84 796
rect 86 792 90 796
rect 92 792 101 796
rect 0 786 4 790
rect 63 786 72 790
rect 74 786 78 790
rect 80 786 84 790
rect 86 786 90 790
rect 92 786 101 790
rect 0 780 4 784
rect 63 780 72 784
rect 74 780 78 784
rect 80 780 84 784
rect 86 780 90 784
rect 92 780 101 784
rect 0 772 4 776
rect 26 772 30 776
rect 32 772 36 776
rect 44 772 48 776
rect 0 766 4 770
rect 14 766 18 770
rect 26 766 30 770
rect 32 766 36 770
rect 44 766 48 770
rect 0 760 4 764
rect 14 760 18 764
rect 26 760 30 764
rect 32 760 36 764
rect 44 760 48 764
rect 0 754 4 758
rect 14 754 18 758
rect 26 754 30 758
rect 32 754 36 758
rect 44 754 48 758
rect 0 748 4 752
rect 14 748 18 752
rect 26 748 30 752
rect 32 748 36 752
rect 44 748 48 752
rect 107 772 111 776
rect 119 772 123 776
rect 107 766 111 770
rect 119 766 123 770
rect 131 766 135 770
rect 107 760 111 764
rect 119 760 123 764
rect 131 760 135 764
rect 107 754 111 758
rect 119 754 123 758
rect 131 754 135 758
rect 107 748 111 752
rect 119 748 123 752
rect 131 748 135 752
rect 0 742 4 746
rect 14 742 18 746
rect 26 742 30 746
rect 32 742 36 746
rect 44 742 48 746
rect 107 742 111 746
rect 119 742 123 746
rect 131 742 135 746
rect 0 736 4 740
rect 14 736 18 740
rect 26 736 30 740
rect 32 736 36 740
rect 44 736 48 740
rect 53 733 57 737
rect 107 736 111 740
rect 119 736 123 740
rect 131 736 135 740
rect 0 723 4 732
rect 53 723 57 727
rect 0 690 4 699
rect 53 695 57 699
rect 0 682 4 686
rect 14 682 18 686
rect 26 682 30 686
rect 32 682 36 686
rect 44 682 48 686
rect 53 685 57 689
rect 107 682 111 686
rect 119 682 123 686
rect 131 682 135 686
rect 0 676 4 680
rect 14 676 18 680
rect 26 676 30 680
rect 32 676 36 680
rect 44 676 48 680
rect 107 676 111 680
rect 119 676 123 680
rect 131 676 135 680
rect 0 670 4 674
rect 14 670 18 674
rect 26 670 30 674
rect 32 670 36 674
rect 44 670 48 674
rect 0 664 4 668
rect 14 664 18 668
rect 26 664 30 668
rect 32 664 36 668
rect 44 664 48 668
rect 0 658 4 662
rect 14 658 18 662
rect 26 658 30 662
rect 32 658 36 662
rect 44 658 48 662
rect 0 652 4 656
rect 14 652 18 656
rect 26 652 30 656
rect 32 652 36 656
rect 44 652 48 656
rect 0 646 4 650
rect 26 646 30 650
rect 32 646 36 650
rect 44 646 48 650
rect 107 670 111 674
rect 119 670 123 674
rect 131 670 135 674
rect 107 664 111 668
rect 119 664 123 668
rect 131 664 135 668
rect 107 658 111 662
rect 119 658 123 662
rect 131 658 135 662
rect 107 652 111 656
rect 119 652 123 656
rect 131 652 135 656
rect 107 646 111 650
rect 119 646 123 650
rect 0 638 4 642
rect 63 638 72 642
rect 74 638 78 642
rect 80 638 84 642
rect 86 638 90 642
rect 92 638 101 642
rect 0 632 4 636
rect 63 632 72 636
rect 74 632 78 636
rect 80 632 84 636
rect 86 632 90 636
rect 92 632 101 636
rect 0 626 4 630
rect 63 626 72 630
rect 74 626 78 630
rect 80 626 84 630
rect 86 626 90 630
rect 92 626 101 630
rect 0 620 4 624
rect 63 620 72 624
rect 74 620 78 624
rect 80 620 84 624
rect 86 620 90 624
rect 92 620 101 624
rect 0 614 4 618
rect 63 614 72 618
rect 74 614 78 618
rect 80 614 84 618
rect 86 614 90 618
rect 92 614 101 618
rect 0 608 4 612
rect 63 608 72 612
rect 74 608 78 612
rect 80 608 84 612
rect 86 608 90 612
rect 92 608 101 612
rect 0 602 4 606
rect 63 602 72 606
rect 74 602 78 606
rect 80 602 84 606
rect 86 602 90 606
rect 92 602 101 606
rect 0 342 4 346
rect 63 342 72 346
rect 74 342 78 346
rect 80 342 84 346
rect 86 342 90 346
rect 92 342 101 346
rect 0 336 4 340
rect 63 336 72 340
rect 74 336 78 340
rect 80 336 84 340
rect 86 336 90 340
rect 92 336 101 340
rect 0 330 4 334
rect 63 330 72 334
rect 74 330 78 334
rect 80 330 84 334
rect 86 330 90 334
rect 92 330 101 334
rect 0 324 4 328
rect 63 324 72 328
rect 74 324 78 328
rect 80 324 84 328
rect 86 324 90 328
rect 92 324 101 328
rect 0 318 4 322
rect 63 318 72 322
rect 74 318 78 322
rect 80 318 84 322
rect 86 318 90 322
rect 92 318 101 322
rect 0 312 4 316
rect 63 312 72 316
rect 74 312 78 316
rect 80 312 84 316
rect 86 312 90 316
rect 92 312 101 316
rect 0 306 4 310
rect 63 306 72 310
rect 74 306 78 310
rect 80 306 84 310
rect 86 306 90 310
rect 92 306 101 310
rect 0 298 4 302
rect 26 298 30 302
rect 32 298 36 302
rect 44 298 48 302
rect 0 292 4 296
rect 14 292 18 296
rect 26 292 30 296
rect 32 292 36 296
rect 44 292 48 296
rect 0 286 4 290
rect 14 286 18 290
rect 26 286 30 290
rect 32 286 36 290
rect 44 286 48 290
rect 0 280 4 284
rect 14 280 18 284
rect 26 280 30 284
rect 32 280 36 284
rect 44 280 48 284
rect 0 274 4 278
rect 14 274 18 278
rect 26 274 30 278
rect 32 274 36 278
rect 44 274 48 278
rect 107 298 111 302
rect 119 298 123 302
rect 107 292 111 296
rect 119 292 123 296
rect 131 292 135 296
rect 107 286 111 290
rect 119 286 123 290
rect 131 286 135 290
rect 107 280 111 284
rect 119 280 123 284
rect 131 280 135 284
rect 107 274 111 278
rect 119 274 123 278
rect 131 274 135 278
rect 0 268 4 272
rect 14 268 18 272
rect 26 268 30 272
rect 32 268 36 272
rect 44 268 48 272
rect 107 268 111 272
rect 119 268 123 272
rect 131 268 135 272
rect 0 262 4 266
rect 14 262 18 266
rect 26 262 30 266
rect 32 262 36 266
rect 44 262 48 266
rect 53 259 57 263
rect 107 262 111 266
rect 119 262 123 266
rect 131 262 135 266
rect 0 249 4 258
rect 53 249 57 253
rect 0 216 4 225
rect 53 221 57 225
rect 0 208 4 212
rect 14 208 18 212
rect 26 208 30 212
rect 32 208 36 212
rect 44 208 48 212
rect 53 211 57 215
rect 107 208 111 212
rect 119 208 123 212
rect 131 208 135 212
rect 0 202 4 206
rect 14 202 18 206
rect 26 202 30 206
rect 32 202 36 206
rect 44 202 48 206
rect 107 202 111 206
rect 119 202 123 206
rect 131 202 135 206
rect 0 196 4 200
rect 14 196 18 200
rect 26 196 30 200
rect 32 196 36 200
rect 44 196 48 200
rect 0 190 4 194
rect 14 190 18 194
rect 26 190 30 194
rect 32 190 36 194
rect 44 190 48 194
rect 0 184 4 188
rect 14 184 18 188
rect 26 184 30 188
rect 32 184 36 188
rect 44 184 48 188
rect 0 178 4 182
rect 14 178 18 182
rect 26 178 30 182
rect 32 178 36 182
rect 44 178 48 182
rect 0 172 4 176
rect 14 172 18 176
rect 26 172 30 176
rect 32 172 36 176
rect 44 172 48 176
rect 107 196 111 200
rect 119 196 123 200
rect 131 196 135 200
rect 107 190 111 194
rect 119 190 123 194
rect 131 190 135 194
rect 107 184 111 188
rect 119 184 123 188
rect 131 184 135 188
rect 107 178 111 182
rect 119 178 123 182
rect 131 178 135 182
rect 107 172 111 176
rect 119 172 123 176
rect 63 164 72 168
rect 74 164 78 168
rect 80 164 84 168
rect 86 164 90 168
rect 92 164 101 168
rect 63 158 72 162
rect 74 158 78 162
rect 80 158 84 162
rect 86 158 90 162
rect 92 158 101 162
rect 63 152 72 156
rect 74 152 78 156
rect 80 152 84 156
rect 86 152 90 156
rect 92 152 101 156
rect 63 146 72 150
rect 74 146 78 150
rect 80 146 84 150
rect 86 146 90 150
rect 92 146 101 150
rect 63 140 72 144
rect 74 140 78 144
rect 80 140 84 144
rect 86 140 90 144
rect 92 140 101 144
rect 63 134 72 138
rect 74 134 78 138
rect 80 134 84 138
rect 86 134 90 138
rect 92 134 101 138
rect 63 128 72 132
rect 74 128 78 132
rect 80 128 84 132
rect 86 128 90 132
rect 92 128 101 132
<< metal2 >>
rect 8 4094 48 4168
rect 4 4090 14 4094
rect 18 4090 26 4094
rect 30 4090 32 4094
rect 36 4090 43 4094
rect 47 4090 48 4094
rect 0 4088 48 4090
rect 4 4084 14 4088
rect 18 4084 26 4088
rect 30 4084 32 4088
rect 36 4084 43 4088
rect 47 4084 48 4088
rect 0 4082 48 4084
rect 4 4078 14 4082
rect 18 4078 26 4082
rect 30 4078 32 4082
rect 36 4078 43 4082
rect 47 4078 48 4082
rect 0 4076 48 4078
rect 4 4072 14 4076
rect 18 4072 26 4076
rect 30 4072 32 4076
rect 36 4072 43 4076
rect 47 4072 48 4076
rect 0 4070 48 4072
rect 4 4066 14 4070
rect 18 4066 26 4070
rect 30 4066 32 4070
rect 36 4066 43 4070
rect 47 4066 48 4070
rect 0 4064 48 4066
rect 4 4060 14 4064
rect 18 4060 26 4064
rect 30 4060 32 4064
rect 36 4060 43 4064
rect 47 4060 48 4064
rect 0 4058 48 4060
rect 4 4054 14 4058
rect 18 4054 26 4058
rect 30 4054 32 4058
rect 36 4054 43 4058
rect 47 4054 48 4058
rect 8 4004 48 4054
rect 4 4000 14 4004
rect 18 4000 26 4004
rect 30 4000 32 4004
rect 36 4000 43 4004
rect 47 4000 48 4004
rect 0 3998 48 4000
rect 4 3994 14 3998
rect 18 3994 26 3998
rect 30 3994 32 3998
rect 36 3994 43 3998
rect 47 3994 48 3998
rect 0 3992 48 3994
rect 4 3988 14 3992
rect 18 3988 26 3992
rect 30 3988 32 3992
rect 36 3988 43 3992
rect 47 3988 48 3992
rect 0 3986 48 3988
rect 4 3982 14 3986
rect 18 3982 26 3986
rect 30 3982 32 3986
rect 36 3982 43 3986
rect 47 3982 48 3986
rect 0 3980 48 3982
rect 4 3976 14 3980
rect 18 3976 26 3980
rect 30 3976 32 3980
rect 36 3976 43 3980
rect 47 3976 48 3980
rect 0 3974 48 3976
rect 4 3970 14 3974
rect 18 3970 26 3974
rect 30 3970 32 3974
rect 36 3970 43 3974
rect 47 3970 48 3974
rect 0 3968 48 3970
rect 4 3964 26 3968
rect 30 3964 32 3968
rect 36 3964 43 3968
rect 47 3964 48 3968
rect 0 3954 4 3956
rect 0 3948 4 3950
rect 0 3942 4 3944
rect 0 3936 4 3938
rect 0 3930 4 3932
rect 0 3924 4 3926
rect 0 3658 4 3660
rect 0 3652 4 3654
rect 0 3646 4 3648
rect 0 3640 4 3642
rect 0 3634 4 3636
rect 0 3628 4 3630
rect 8 3620 48 3964
rect 4 3616 26 3620
rect 30 3616 32 3620
rect 36 3616 44 3620
rect 0 3614 48 3616
rect 4 3610 14 3614
rect 18 3610 26 3614
rect 30 3610 32 3614
rect 36 3610 44 3614
rect 0 3608 48 3610
rect 4 3604 14 3608
rect 18 3604 26 3608
rect 30 3604 32 3608
rect 36 3604 44 3608
rect 0 3602 48 3604
rect 4 3598 14 3602
rect 18 3598 26 3602
rect 30 3598 32 3602
rect 36 3598 44 3602
rect 0 3596 48 3598
rect 4 3592 14 3596
rect 18 3592 26 3596
rect 30 3592 32 3596
rect 36 3592 44 3596
rect 0 3590 48 3592
rect 4 3586 14 3590
rect 18 3586 26 3590
rect 30 3586 32 3590
rect 36 3586 44 3590
rect 0 3584 48 3586
rect 4 3580 14 3584
rect 18 3580 26 3584
rect 30 3580 32 3584
rect 36 3580 44 3584
rect 8 3530 48 3580
rect 4 3526 14 3530
rect 18 3526 26 3530
rect 30 3526 32 3530
rect 36 3526 44 3530
rect 0 3524 48 3526
rect 4 3520 14 3524
rect 18 3520 26 3524
rect 30 3520 32 3524
rect 36 3520 44 3524
rect 0 3518 48 3520
rect 4 3514 14 3518
rect 18 3514 26 3518
rect 30 3514 32 3518
rect 36 3514 44 3518
rect 0 3512 48 3514
rect 4 3508 14 3512
rect 18 3508 26 3512
rect 30 3508 32 3512
rect 36 3508 44 3512
rect 0 3506 48 3508
rect 4 3502 14 3506
rect 18 3502 26 3506
rect 30 3502 32 3506
rect 36 3502 44 3506
rect 0 3500 48 3502
rect 4 3496 14 3500
rect 18 3496 26 3500
rect 30 3496 32 3500
rect 36 3496 44 3500
rect 0 3494 48 3496
rect 4 3490 26 3494
rect 30 3490 32 3494
rect 36 3490 44 3494
rect 0 3480 4 3482
rect 0 3474 4 3476
rect 0 3468 4 3470
rect 0 3462 4 3464
rect 0 3456 4 3458
rect 0 3450 4 3452
rect 0 3184 4 3186
rect 0 3178 4 3180
rect 0 3172 4 3174
rect 0 3166 4 3168
rect 0 3160 4 3162
rect 0 3154 4 3156
rect 8 3146 48 3490
rect 4 3142 26 3146
rect 30 3142 32 3146
rect 36 3142 44 3146
rect 0 3140 48 3142
rect 4 3136 14 3140
rect 18 3136 26 3140
rect 30 3136 32 3140
rect 36 3136 44 3140
rect 0 3134 48 3136
rect 4 3130 14 3134
rect 18 3130 26 3134
rect 30 3130 32 3134
rect 36 3130 44 3134
rect 0 3128 48 3130
rect 4 3124 14 3128
rect 18 3124 26 3128
rect 30 3124 32 3128
rect 36 3124 44 3128
rect 0 3122 48 3124
rect 4 3118 14 3122
rect 18 3118 26 3122
rect 30 3118 32 3122
rect 36 3118 44 3122
rect 0 3116 48 3118
rect 4 3112 14 3116
rect 18 3112 26 3116
rect 30 3112 32 3116
rect 36 3112 44 3116
rect 0 3110 48 3112
rect 4 3106 14 3110
rect 18 3106 26 3110
rect 30 3106 32 3110
rect 36 3106 44 3110
rect 8 3056 48 3106
rect 4 3052 14 3056
rect 18 3052 26 3056
rect 30 3052 32 3056
rect 36 3052 44 3056
rect 0 3050 48 3052
rect 4 3046 14 3050
rect 18 3046 26 3050
rect 30 3046 32 3050
rect 36 3046 44 3050
rect 0 3044 48 3046
rect 4 3040 14 3044
rect 18 3040 26 3044
rect 30 3040 32 3044
rect 36 3040 44 3044
rect 0 3038 48 3040
rect 4 3034 14 3038
rect 18 3034 26 3038
rect 30 3034 32 3038
rect 36 3034 44 3038
rect 0 3032 48 3034
rect 4 3028 14 3032
rect 18 3028 26 3032
rect 30 3028 32 3032
rect 36 3028 44 3032
rect 0 3026 48 3028
rect 4 3022 14 3026
rect 18 3022 26 3026
rect 30 3022 32 3026
rect 36 3022 44 3026
rect 0 3020 48 3022
rect 4 3016 26 3020
rect 30 3016 32 3020
rect 36 3016 44 3020
rect 0 3006 4 3008
rect 0 3000 4 3002
rect 0 2994 4 2996
rect 0 2988 4 2990
rect 0 2982 4 2984
rect 0 2976 4 2978
rect 0 2710 4 2712
rect 0 2704 4 2706
rect 0 2698 4 2700
rect 0 2692 4 2694
rect 0 2686 4 2688
rect 0 2680 4 2682
rect 8 2672 48 3016
rect 4 2668 26 2672
rect 30 2668 32 2672
rect 36 2668 44 2672
rect 0 2666 48 2668
rect 4 2662 14 2666
rect 18 2662 26 2666
rect 30 2662 32 2666
rect 36 2662 44 2666
rect 0 2660 48 2662
rect 4 2656 14 2660
rect 18 2656 26 2660
rect 30 2656 32 2660
rect 36 2656 44 2660
rect 0 2654 48 2656
rect 4 2650 14 2654
rect 18 2650 26 2654
rect 30 2650 32 2654
rect 36 2650 44 2654
rect 0 2648 48 2650
rect 4 2644 14 2648
rect 18 2644 26 2648
rect 30 2644 32 2648
rect 36 2644 44 2648
rect 0 2642 48 2644
rect 4 2638 14 2642
rect 18 2638 26 2642
rect 30 2638 32 2642
rect 36 2638 44 2642
rect 0 2636 48 2638
rect 4 2632 14 2636
rect 18 2632 26 2636
rect 30 2632 32 2636
rect 36 2632 44 2636
rect 8 2582 48 2632
rect 4 2578 14 2582
rect 18 2578 26 2582
rect 30 2578 32 2582
rect 36 2578 44 2582
rect 0 2576 48 2578
rect 4 2572 14 2576
rect 18 2572 26 2576
rect 30 2572 32 2576
rect 36 2572 44 2576
rect 0 2570 48 2572
rect 4 2566 14 2570
rect 18 2566 26 2570
rect 30 2566 32 2570
rect 36 2566 44 2570
rect 0 2564 48 2566
rect 4 2560 14 2564
rect 18 2560 26 2564
rect 30 2560 32 2564
rect 36 2560 44 2564
rect 0 2558 48 2560
rect 4 2554 14 2558
rect 18 2554 26 2558
rect 30 2554 32 2558
rect 36 2554 44 2558
rect 0 2552 48 2554
rect 4 2548 14 2552
rect 18 2548 26 2552
rect 30 2548 32 2552
rect 36 2548 44 2552
rect 0 2546 48 2548
rect 4 2542 26 2546
rect 30 2542 32 2546
rect 36 2542 44 2546
rect 0 2532 4 2534
rect 0 2526 4 2528
rect 0 2520 4 2522
rect 0 2514 4 2516
rect 0 2508 4 2510
rect 0 2502 4 2504
rect 0 2236 4 2238
rect 0 2230 4 2232
rect 0 2224 4 2226
rect 0 2218 4 2220
rect 0 2212 4 2214
rect 0 2206 4 2208
rect 8 2198 48 2542
rect 4 2194 26 2198
rect 30 2194 32 2198
rect 36 2194 44 2198
rect 0 2192 48 2194
rect 4 2188 14 2192
rect 18 2188 26 2192
rect 30 2188 32 2192
rect 36 2188 44 2192
rect 0 2186 48 2188
rect 4 2182 14 2186
rect 18 2182 26 2186
rect 30 2182 32 2186
rect 36 2182 44 2186
rect 0 2180 48 2182
rect 4 2176 14 2180
rect 18 2176 26 2180
rect 30 2176 32 2180
rect 36 2176 44 2180
rect 0 2174 48 2176
rect 4 2170 14 2174
rect 18 2170 26 2174
rect 30 2170 32 2174
rect 36 2170 44 2174
rect 0 2168 48 2170
rect 4 2164 14 2168
rect 18 2164 26 2168
rect 30 2164 32 2168
rect 36 2164 44 2168
rect 0 2162 48 2164
rect 4 2158 14 2162
rect 18 2158 26 2162
rect 30 2158 32 2162
rect 36 2158 44 2162
rect 8 2108 48 2158
rect 4 2104 14 2108
rect 18 2104 26 2108
rect 30 2104 32 2108
rect 36 2104 44 2108
rect 0 2102 48 2104
rect 4 2098 14 2102
rect 18 2098 26 2102
rect 30 2098 32 2102
rect 36 2098 44 2102
rect 0 2096 48 2098
rect 4 2092 14 2096
rect 18 2092 26 2096
rect 30 2092 32 2096
rect 36 2092 44 2096
rect 0 2090 48 2092
rect 4 2086 14 2090
rect 18 2086 26 2090
rect 30 2086 32 2090
rect 36 2086 44 2090
rect 0 2084 48 2086
rect 4 2080 14 2084
rect 18 2080 26 2084
rect 30 2080 32 2084
rect 36 2080 44 2084
rect 0 2078 48 2080
rect 4 2074 14 2078
rect 18 2074 26 2078
rect 30 2074 32 2078
rect 36 2074 44 2078
rect 0 2072 48 2074
rect 4 2068 26 2072
rect 30 2068 32 2072
rect 36 2068 44 2072
rect 0 2058 4 2060
rect 0 2052 4 2054
rect 0 2046 4 2048
rect 0 2040 4 2042
rect 0 2034 4 2036
rect 0 2028 4 2030
rect 0 1762 4 1764
rect 0 1756 4 1758
rect 0 1750 4 1752
rect 0 1744 4 1746
rect 0 1738 4 1740
rect 0 1732 4 1734
rect 8 1724 48 2068
rect 4 1720 26 1724
rect 30 1720 32 1724
rect 36 1720 44 1724
rect 0 1718 48 1720
rect 4 1714 14 1718
rect 18 1714 26 1718
rect 30 1714 32 1718
rect 36 1714 44 1718
rect 0 1712 48 1714
rect 4 1708 14 1712
rect 18 1708 26 1712
rect 30 1708 32 1712
rect 36 1708 44 1712
rect 0 1706 48 1708
rect 4 1702 14 1706
rect 18 1702 26 1706
rect 30 1702 32 1706
rect 36 1702 44 1706
rect 0 1700 48 1702
rect 4 1696 14 1700
rect 18 1696 26 1700
rect 30 1696 32 1700
rect 36 1696 44 1700
rect 0 1694 48 1696
rect 4 1690 14 1694
rect 18 1690 26 1694
rect 30 1690 32 1694
rect 36 1690 44 1694
rect 0 1688 48 1690
rect 4 1684 14 1688
rect 18 1684 26 1688
rect 30 1684 32 1688
rect 36 1684 44 1688
rect 8 1634 48 1684
rect 4 1630 14 1634
rect 18 1630 26 1634
rect 30 1630 32 1634
rect 36 1630 44 1634
rect 0 1628 48 1630
rect 4 1624 14 1628
rect 18 1624 26 1628
rect 30 1624 32 1628
rect 36 1624 44 1628
rect 0 1622 48 1624
rect 4 1618 14 1622
rect 18 1618 26 1622
rect 30 1618 32 1622
rect 36 1618 44 1622
rect 0 1616 48 1618
rect 4 1612 14 1616
rect 18 1612 26 1616
rect 30 1612 32 1616
rect 36 1612 44 1616
rect 0 1610 48 1612
rect 4 1606 14 1610
rect 18 1606 26 1610
rect 30 1606 32 1610
rect 36 1606 44 1610
rect 0 1604 48 1606
rect 4 1600 14 1604
rect 18 1600 26 1604
rect 30 1600 32 1604
rect 36 1600 44 1604
rect 0 1598 48 1600
rect 4 1594 26 1598
rect 30 1594 32 1598
rect 36 1594 44 1598
rect 0 1584 4 1586
rect 0 1578 4 1580
rect 0 1572 4 1574
rect 0 1566 4 1568
rect 0 1560 4 1562
rect 0 1554 4 1556
rect 0 1288 4 1290
rect 0 1282 4 1284
rect 0 1276 4 1278
rect 0 1270 4 1272
rect 0 1264 4 1266
rect 0 1258 4 1260
rect 8 1250 48 1594
rect 4 1246 26 1250
rect 30 1246 32 1250
rect 36 1246 44 1250
rect 0 1244 48 1246
rect 4 1240 14 1244
rect 18 1240 26 1244
rect 30 1240 32 1244
rect 36 1240 44 1244
rect 0 1238 48 1240
rect 4 1234 14 1238
rect 18 1234 26 1238
rect 30 1234 32 1238
rect 36 1234 44 1238
rect 0 1232 48 1234
rect 4 1228 14 1232
rect 18 1228 26 1232
rect 30 1228 32 1232
rect 36 1228 44 1232
rect 0 1226 48 1228
rect 4 1222 14 1226
rect 18 1222 26 1226
rect 30 1222 32 1226
rect 36 1222 44 1226
rect 0 1220 48 1222
rect 4 1216 14 1220
rect 18 1216 26 1220
rect 30 1216 32 1220
rect 36 1216 44 1220
rect 0 1214 48 1216
rect 4 1210 14 1214
rect 18 1210 26 1214
rect 30 1210 32 1214
rect 36 1210 44 1214
rect 8 1160 48 1210
rect 4 1156 14 1160
rect 18 1156 26 1160
rect 30 1156 32 1160
rect 36 1156 44 1160
rect 0 1154 48 1156
rect 4 1150 14 1154
rect 18 1150 26 1154
rect 30 1150 32 1154
rect 36 1150 44 1154
rect 0 1148 48 1150
rect 4 1144 14 1148
rect 18 1144 26 1148
rect 30 1144 32 1148
rect 36 1144 44 1148
rect 0 1142 48 1144
rect 4 1138 14 1142
rect 18 1138 26 1142
rect 30 1138 32 1142
rect 36 1138 44 1142
rect 0 1136 48 1138
rect 4 1132 14 1136
rect 18 1132 26 1136
rect 30 1132 32 1136
rect 36 1132 44 1136
rect 0 1130 48 1132
rect 4 1126 14 1130
rect 18 1126 26 1130
rect 30 1126 32 1130
rect 36 1126 44 1130
rect 0 1124 48 1126
rect 4 1120 26 1124
rect 30 1120 32 1124
rect 36 1120 44 1124
rect 0 1110 4 1112
rect 0 1104 4 1106
rect 0 1098 4 1100
rect 0 1092 4 1094
rect 0 1086 4 1088
rect 0 1080 4 1082
rect 0 814 4 816
rect 0 808 4 810
rect 0 802 4 804
rect 0 796 4 798
rect 0 790 4 792
rect 0 784 4 786
rect 8 776 48 1120
rect 4 772 26 776
rect 30 772 32 776
rect 36 772 44 776
rect 0 770 48 772
rect 4 766 14 770
rect 18 766 26 770
rect 30 766 32 770
rect 36 766 44 770
rect 0 764 48 766
rect 4 760 14 764
rect 18 760 26 764
rect 30 760 32 764
rect 36 760 44 764
rect 0 758 48 760
rect 4 754 14 758
rect 18 754 26 758
rect 30 754 32 758
rect 36 754 44 758
rect 0 752 48 754
rect 4 748 14 752
rect 18 748 26 752
rect 30 748 32 752
rect 36 748 44 752
rect 0 746 48 748
rect 4 742 14 746
rect 18 742 26 746
rect 30 742 32 746
rect 36 742 44 746
rect 0 740 48 742
rect 4 736 14 740
rect 18 736 26 740
rect 30 736 32 740
rect 36 736 44 740
rect 8 686 48 736
rect 4 682 14 686
rect 18 682 26 686
rect 30 682 32 686
rect 36 682 44 686
rect 0 680 48 682
rect 4 676 14 680
rect 18 676 26 680
rect 30 676 32 680
rect 36 676 44 680
rect 0 674 48 676
rect 4 670 14 674
rect 18 670 26 674
rect 30 670 32 674
rect 36 670 44 674
rect 0 668 48 670
rect 4 664 14 668
rect 18 664 26 668
rect 30 664 32 668
rect 36 664 44 668
rect 0 662 48 664
rect 4 658 14 662
rect 18 658 26 662
rect 30 658 32 662
rect 36 658 44 662
rect 0 656 48 658
rect 4 652 14 656
rect 18 652 26 656
rect 30 652 32 656
rect 36 652 44 656
rect 0 650 48 652
rect 4 646 26 650
rect 30 646 32 650
rect 36 646 44 650
rect 0 636 4 638
rect 0 630 4 632
rect 0 624 4 626
rect 0 618 4 620
rect 0 612 4 614
rect 0 606 4 608
rect 0 340 4 342
rect 0 334 4 336
rect 0 328 4 330
rect 0 322 4 324
rect 0 316 4 318
rect 0 310 4 312
rect 8 302 48 646
rect 4 298 26 302
rect 30 298 32 302
rect 36 298 44 302
rect 0 296 48 298
rect 4 292 14 296
rect 18 292 26 296
rect 30 292 32 296
rect 36 292 44 296
rect 0 290 48 292
rect 4 286 14 290
rect 18 286 26 290
rect 30 286 32 290
rect 36 286 44 290
rect 0 284 48 286
rect 4 280 14 284
rect 18 280 26 284
rect 30 280 32 284
rect 36 280 44 284
rect 0 278 48 280
rect 4 274 14 278
rect 18 274 26 278
rect 30 274 32 278
rect 36 274 44 278
rect 0 272 48 274
rect 4 268 14 272
rect 18 268 26 272
rect 30 268 32 272
rect 36 268 44 272
rect 0 266 48 268
rect 4 262 14 266
rect 18 262 26 266
rect 30 262 32 266
rect 36 262 44 266
rect 8 212 48 262
rect 4 208 14 212
rect 18 208 26 212
rect 30 208 32 212
rect 36 208 44 212
rect 0 206 48 208
rect 4 202 14 206
rect 18 202 26 206
rect 30 202 32 206
rect 36 202 44 206
rect 0 200 48 202
rect 4 196 14 200
rect 18 196 26 200
rect 30 196 32 200
rect 36 196 44 200
rect 0 194 48 196
rect 4 190 14 194
rect 18 190 26 194
rect 30 190 32 194
rect 36 190 44 194
rect 0 188 48 190
rect 4 184 14 188
rect 18 184 26 188
rect 30 184 32 188
rect 36 184 44 188
rect 0 182 48 184
rect 4 178 14 182
rect 18 178 26 182
rect 30 178 32 182
rect 36 178 44 182
rect 0 176 48 178
rect 4 172 14 176
rect 18 172 26 176
rect 30 172 32 176
rect 36 172 44 176
rect 8 98 48 172
rect 52 4055 58 4172
rect 52 4051 53 4055
rect 57 4051 58 4055
rect 52 4045 58 4051
rect 52 4041 53 4045
rect 57 4041 58 4045
rect 52 4017 58 4041
rect 52 4013 53 4017
rect 57 4013 58 4017
rect 52 4007 58 4013
rect 52 4003 53 4007
rect 57 4003 58 4007
rect 52 3581 58 4003
rect 52 3577 53 3581
rect 57 3577 58 3581
rect 52 3571 58 3577
rect 52 3567 53 3571
rect 57 3567 58 3571
rect 52 3543 58 3567
rect 52 3539 53 3543
rect 57 3539 58 3543
rect 52 3533 58 3539
rect 52 3529 53 3533
rect 57 3529 58 3533
rect 52 3107 58 3529
rect 52 3103 53 3107
rect 57 3103 58 3107
rect 52 3097 58 3103
rect 52 3093 53 3097
rect 57 3093 58 3097
rect 52 3069 58 3093
rect 52 3065 53 3069
rect 57 3065 58 3069
rect 52 3059 58 3065
rect 52 3055 53 3059
rect 57 3055 58 3059
rect 52 2633 58 3055
rect 52 2629 53 2633
rect 57 2629 58 2633
rect 52 2623 58 2629
rect 52 2619 53 2623
rect 57 2619 58 2623
rect 52 2595 58 2619
rect 52 2591 53 2595
rect 57 2591 58 2595
rect 52 2585 58 2591
rect 52 2581 53 2585
rect 57 2581 58 2585
rect 52 2159 58 2581
rect 52 2155 53 2159
rect 57 2155 58 2159
rect 52 2149 58 2155
rect 52 2145 53 2149
rect 57 2145 58 2149
rect 52 2121 58 2145
rect 52 2117 53 2121
rect 57 2117 58 2121
rect 52 2111 58 2117
rect 52 2107 53 2111
rect 57 2107 58 2111
rect 52 1685 58 2107
rect 52 1681 53 1685
rect 57 1681 58 1685
rect 52 1675 58 1681
rect 52 1671 53 1675
rect 57 1671 58 1675
rect 52 1647 58 1671
rect 52 1643 53 1647
rect 57 1643 58 1647
rect 52 1637 58 1643
rect 52 1633 53 1637
rect 57 1633 58 1637
rect 52 1211 58 1633
rect 52 1207 53 1211
rect 57 1207 58 1211
rect 52 1201 58 1207
rect 52 1197 53 1201
rect 57 1197 58 1201
rect 52 1173 58 1197
rect 52 1169 53 1173
rect 57 1169 58 1173
rect 52 1163 58 1169
rect 52 1159 53 1163
rect 57 1159 58 1163
rect 52 737 58 1159
rect 52 733 53 737
rect 57 733 58 737
rect 52 727 58 733
rect 52 723 53 727
rect 57 723 58 727
rect 52 699 58 723
rect 52 695 53 699
rect 57 695 58 699
rect 52 689 58 695
rect 52 685 53 689
rect 57 685 58 689
rect 52 263 58 685
rect 52 259 53 263
rect 57 259 58 263
rect 52 253 58 259
rect 52 249 53 253
rect 57 249 58 253
rect 52 225 58 249
rect 52 221 53 225
rect 57 221 58 225
rect 52 215 58 221
rect 52 211 53 215
rect 57 211 58 215
rect 52 94 58 211
rect 62 4138 102 4182
rect 62 4134 63 4138
rect 72 4134 74 4138
rect 78 4134 80 4138
rect 84 4134 86 4138
rect 90 4134 92 4138
rect 101 4134 102 4138
rect 62 4132 102 4134
rect 62 4128 63 4132
rect 72 4128 74 4132
rect 78 4128 80 4132
rect 84 4128 86 4132
rect 90 4128 92 4132
rect 101 4128 102 4132
rect 62 4126 102 4128
rect 62 4122 63 4126
rect 72 4122 74 4126
rect 78 4122 80 4126
rect 84 4122 86 4126
rect 90 4122 92 4126
rect 101 4122 102 4126
rect 62 4120 102 4122
rect 62 4116 63 4120
rect 72 4116 74 4120
rect 78 4116 80 4120
rect 84 4116 86 4120
rect 90 4116 92 4120
rect 101 4116 102 4120
rect 62 4114 102 4116
rect 62 4110 63 4114
rect 72 4110 74 4114
rect 78 4110 80 4114
rect 84 4110 86 4114
rect 90 4110 92 4114
rect 101 4110 102 4114
rect 62 4108 102 4110
rect 62 4104 63 4108
rect 72 4104 74 4108
rect 78 4104 80 4108
rect 84 4104 86 4108
rect 90 4104 92 4108
rect 101 4104 102 4108
rect 62 4102 102 4104
rect 62 4098 63 4102
rect 72 4098 74 4102
rect 78 4098 80 4102
rect 84 4098 86 4102
rect 90 4098 92 4102
rect 101 4098 102 4102
rect 62 3960 102 4098
rect 62 3956 63 3960
rect 72 3956 74 3960
rect 78 3956 80 3960
rect 84 3956 86 3960
rect 90 3956 92 3960
rect 101 3956 102 3960
rect 62 3954 102 3956
rect 62 3950 63 3954
rect 72 3950 74 3954
rect 78 3950 80 3954
rect 84 3950 86 3954
rect 90 3950 92 3954
rect 101 3950 102 3954
rect 62 3948 102 3950
rect 62 3944 63 3948
rect 72 3944 74 3948
rect 78 3944 80 3948
rect 84 3944 86 3948
rect 90 3944 92 3948
rect 101 3944 102 3948
rect 62 3942 102 3944
rect 62 3938 63 3942
rect 72 3938 74 3942
rect 78 3938 80 3942
rect 84 3938 86 3942
rect 90 3938 92 3942
rect 101 3938 102 3942
rect 62 3936 102 3938
rect 62 3932 63 3936
rect 72 3932 74 3936
rect 78 3932 80 3936
rect 84 3932 86 3936
rect 90 3932 92 3936
rect 101 3932 102 3936
rect 62 3930 102 3932
rect 62 3926 63 3930
rect 72 3926 74 3930
rect 78 3926 80 3930
rect 84 3926 86 3930
rect 90 3926 92 3930
rect 101 3926 102 3930
rect 62 3924 102 3926
rect 62 3920 63 3924
rect 72 3920 74 3924
rect 78 3920 80 3924
rect 84 3920 86 3924
rect 90 3920 92 3924
rect 101 3920 102 3924
rect 62 3664 102 3920
rect 62 3660 63 3664
rect 72 3660 74 3664
rect 78 3660 80 3664
rect 84 3660 86 3664
rect 90 3660 92 3664
rect 101 3660 102 3664
rect 62 3658 102 3660
rect 62 3654 63 3658
rect 72 3654 74 3658
rect 78 3654 80 3658
rect 84 3654 86 3658
rect 90 3654 92 3658
rect 101 3654 102 3658
rect 62 3652 102 3654
rect 62 3648 63 3652
rect 72 3648 74 3652
rect 78 3648 80 3652
rect 84 3648 86 3652
rect 90 3648 92 3652
rect 101 3648 102 3652
rect 62 3646 102 3648
rect 62 3642 63 3646
rect 72 3642 74 3646
rect 78 3642 80 3646
rect 84 3642 86 3646
rect 90 3642 92 3646
rect 101 3642 102 3646
rect 62 3640 102 3642
rect 62 3636 63 3640
rect 72 3636 74 3640
rect 78 3636 80 3640
rect 84 3636 86 3640
rect 90 3636 92 3640
rect 101 3636 102 3640
rect 62 3634 102 3636
rect 62 3630 63 3634
rect 72 3630 74 3634
rect 78 3630 80 3634
rect 84 3630 86 3634
rect 90 3630 92 3634
rect 101 3630 102 3634
rect 62 3628 102 3630
rect 62 3624 63 3628
rect 72 3624 74 3628
rect 78 3624 80 3628
rect 84 3624 86 3628
rect 90 3624 92 3628
rect 101 3624 102 3628
rect 62 3486 102 3624
rect 62 3482 63 3486
rect 72 3482 74 3486
rect 78 3482 80 3486
rect 84 3482 86 3486
rect 90 3482 92 3486
rect 101 3482 102 3486
rect 62 3480 102 3482
rect 62 3476 63 3480
rect 72 3476 74 3480
rect 78 3476 80 3480
rect 84 3476 86 3480
rect 90 3476 92 3480
rect 101 3476 102 3480
rect 62 3474 102 3476
rect 62 3470 63 3474
rect 72 3470 74 3474
rect 78 3470 80 3474
rect 84 3470 86 3474
rect 90 3470 92 3474
rect 101 3470 102 3474
rect 62 3468 102 3470
rect 62 3464 63 3468
rect 72 3464 74 3468
rect 78 3464 80 3468
rect 84 3464 86 3468
rect 90 3464 92 3468
rect 101 3464 102 3468
rect 62 3462 102 3464
rect 62 3458 63 3462
rect 72 3458 74 3462
rect 78 3458 80 3462
rect 84 3458 86 3462
rect 90 3458 92 3462
rect 101 3458 102 3462
rect 62 3456 102 3458
rect 62 3452 63 3456
rect 72 3452 74 3456
rect 78 3452 80 3456
rect 84 3452 86 3456
rect 90 3452 92 3456
rect 101 3452 102 3456
rect 62 3450 102 3452
rect 62 3446 63 3450
rect 72 3446 74 3450
rect 78 3446 80 3450
rect 84 3446 86 3450
rect 90 3446 92 3450
rect 101 3446 102 3450
rect 62 3190 102 3446
rect 62 3186 63 3190
rect 72 3186 74 3190
rect 78 3186 80 3190
rect 84 3186 86 3190
rect 90 3186 92 3190
rect 101 3186 102 3190
rect 62 3184 102 3186
rect 62 3180 63 3184
rect 72 3180 74 3184
rect 78 3180 80 3184
rect 84 3180 86 3184
rect 90 3180 92 3184
rect 101 3180 102 3184
rect 62 3178 102 3180
rect 62 3174 63 3178
rect 72 3174 74 3178
rect 78 3174 80 3178
rect 84 3174 86 3178
rect 90 3174 92 3178
rect 101 3174 102 3178
rect 62 3172 102 3174
rect 62 3168 63 3172
rect 72 3168 74 3172
rect 78 3168 80 3172
rect 84 3168 86 3172
rect 90 3168 92 3172
rect 101 3168 102 3172
rect 62 3166 102 3168
rect 62 3162 63 3166
rect 72 3162 74 3166
rect 78 3162 80 3166
rect 84 3162 86 3166
rect 90 3162 92 3166
rect 101 3162 102 3166
rect 62 3160 102 3162
rect 62 3156 63 3160
rect 72 3156 74 3160
rect 78 3156 80 3160
rect 84 3156 86 3160
rect 90 3156 92 3160
rect 101 3156 102 3160
rect 62 3154 102 3156
rect 62 3150 63 3154
rect 72 3150 74 3154
rect 78 3150 80 3154
rect 84 3150 86 3154
rect 90 3150 92 3154
rect 101 3150 102 3154
rect 62 3012 102 3150
rect 62 3008 63 3012
rect 72 3008 74 3012
rect 78 3008 80 3012
rect 84 3008 86 3012
rect 90 3008 92 3012
rect 101 3008 102 3012
rect 62 3006 102 3008
rect 62 3002 63 3006
rect 72 3002 74 3006
rect 78 3002 80 3006
rect 84 3002 86 3006
rect 90 3002 92 3006
rect 101 3002 102 3006
rect 62 3000 102 3002
rect 62 2996 63 3000
rect 72 2996 74 3000
rect 78 2996 80 3000
rect 84 2996 86 3000
rect 90 2996 92 3000
rect 101 2996 102 3000
rect 62 2994 102 2996
rect 62 2990 63 2994
rect 72 2990 74 2994
rect 78 2990 80 2994
rect 84 2990 86 2994
rect 90 2990 92 2994
rect 101 2990 102 2994
rect 62 2988 102 2990
rect 62 2984 63 2988
rect 72 2984 74 2988
rect 78 2984 80 2988
rect 84 2984 86 2988
rect 90 2984 92 2988
rect 101 2984 102 2988
rect 62 2982 102 2984
rect 62 2978 63 2982
rect 72 2978 74 2982
rect 78 2978 80 2982
rect 84 2978 86 2982
rect 90 2978 92 2982
rect 101 2978 102 2982
rect 62 2976 102 2978
rect 62 2972 63 2976
rect 72 2972 74 2976
rect 78 2972 80 2976
rect 84 2972 86 2976
rect 90 2972 92 2976
rect 101 2972 102 2976
rect 62 2716 102 2972
rect 62 2712 63 2716
rect 72 2712 74 2716
rect 78 2712 80 2716
rect 84 2712 86 2716
rect 90 2712 92 2716
rect 101 2712 102 2716
rect 62 2710 102 2712
rect 62 2706 63 2710
rect 72 2706 74 2710
rect 78 2706 80 2710
rect 84 2706 86 2710
rect 90 2706 92 2710
rect 101 2706 102 2710
rect 62 2704 102 2706
rect 62 2700 63 2704
rect 72 2700 74 2704
rect 78 2700 80 2704
rect 84 2700 86 2704
rect 90 2700 92 2704
rect 101 2700 102 2704
rect 62 2698 102 2700
rect 62 2694 63 2698
rect 72 2694 74 2698
rect 78 2694 80 2698
rect 84 2694 86 2698
rect 90 2694 92 2698
rect 101 2694 102 2698
rect 62 2692 102 2694
rect 62 2688 63 2692
rect 72 2688 74 2692
rect 78 2688 80 2692
rect 84 2688 86 2692
rect 90 2688 92 2692
rect 101 2688 102 2692
rect 62 2686 102 2688
rect 62 2682 63 2686
rect 72 2682 74 2686
rect 78 2682 80 2686
rect 84 2682 86 2686
rect 90 2682 92 2686
rect 101 2682 102 2686
rect 62 2680 102 2682
rect 62 2676 63 2680
rect 72 2676 74 2680
rect 78 2676 80 2680
rect 84 2676 86 2680
rect 90 2676 92 2680
rect 101 2676 102 2680
rect 62 2538 102 2676
rect 62 2534 63 2538
rect 72 2534 74 2538
rect 78 2534 80 2538
rect 84 2534 86 2538
rect 90 2534 92 2538
rect 101 2534 102 2538
rect 62 2532 102 2534
rect 62 2528 63 2532
rect 72 2528 74 2532
rect 78 2528 80 2532
rect 84 2528 86 2532
rect 90 2528 92 2532
rect 101 2528 102 2532
rect 62 2526 102 2528
rect 62 2522 63 2526
rect 72 2522 74 2526
rect 78 2522 80 2526
rect 84 2522 86 2526
rect 90 2522 92 2526
rect 101 2522 102 2526
rect 62 2520 102 2522
rect 62 2516 63 2520
rect 72 2516 74 2520
rect 78 2516 80 2520
rect 84 2516 86 2520
rect 90 2516 92 2520
rect 101 2516 102 2520
rect 62 2514 102 2516
rect 62 2510 63 2514
rect 72 2510 74 2514
rect 78 2510 80 2514
rect 84 2510 86 2514
rect 90 2510 92 2514
rect 101 2510 102 2514
rect 62 2508 102 2510
rect 62 2504 63 2508
rect 72 2504 74 2508
rect 78 2504 80 2508
rect 84 2504 86 2508
rect 90 2504 92 2508
rect 101 2504 102 2508
rect 62 2502 102 2504
rect 62 2498 63 2502
rect 72 2498 74 2502
rect 78 2498 80 2502
rect 84 2498 86 2502
rect 90 2498 92 2502
rect 101 2498 102 2502
rect 62 2242 102 2498
rect 62 2238 63 2242
rect 72 2238 74 2242
rect 78 2238 80 2242
rect 84 2238 86 2242
rect 90 2238 92 2242
rect 101 2238 102 2242
rect 62 2236 102 2238
rect 62 2232 63 2236
rect 72 2232 74 2236
rect 78 2232 80 2236
rect 84 2232 86 2236
rect 90 2232 92 2236
rect 101 2232 102 2236
rect 62 2230 102 2232
rect 62 2226 63 2230
rect 72 2226 74 2230
rect 78 2226 80 2230
rect 84 2226 86 2230
rect 90 2226 92 2230
rect 101 2226 102 2230
rect 62 2224 102 2226
rect 62 2220 63 2224
rect 72 2220 74 2224
rect 78 2220 80 2224
rect 84 2220 86 2224
rect 90 2220 92 2224
rect 101 2220 102 2224
rect 62 2218 102 2220
rect 62 2214 63 2218
rect 72 2214 74 2218
rect 78 2214 80 2218
rect 84 2214 86 2218
rect 90 2214 92 2218
rect 101 2214 102 2218
rect 62 2212 102 2214
rect 62 2208 63 2212
rect 72 2208 74 2212
rect 78 2208 80 2212
rect 84 2208 86 2212
rect 90 2208 92 2212
rect 101 2208 102 2212
rect 62 2206 102 2208
rect 62 2202 63 2206
rect 72 2202 74 2206
rect 78 2202 80 2206
rect 84 2202 86 2206
rect 90 2202 92 2206
rect 101 2202 102 2206
rect 62 2064 102 2202
rect 62 2060 63 2064
rect 72 2060 74 2064
rect 78 2060 80 2064
rect 84 2060 86 2064
rect 90 2060 92 2064
rect 101 2060 102 2064
rect 62 2058 102 2060
rect 62 2054 63 2058
rect 72 2054 74 2058
rect 78 2054 80 2058
rect 84 2054 86 2058
rect 90 2054 92 2058
rect 101 2054 102 2058
rect 62 2052 102 2054
rect 62 2048 63 2052
rect 72 2048 74 2052
rect 78 2048 80 2052
rect 84 2048 86 2052
rect 90 2048 92 2052
rect 101 2048 102 2052
rect 62 2046 102 2048
rect 62 2042 63 2046
rect 72 2042 74 2046
rect 78 2042 80 2046
rect 84 2042 86 2046
rect 90 2042 92 2046
rect 101 2042 102 2046
rect 62 2040 102 2042
rect 62 2036 63 2040
rect 72 2036 74 2040
rect 78 2036 80 2040
rect 84 2036 86 2040
rect 90 2036 92 2040
rect 101 2036 102 2040
rect 62 2034 102 2036
rect 62 2030 63 2034
rect 72 2030 74 2034
rect 78 2030 80 2034
rect 84 2030 86 2034
rect 90 2030 92 2034
rect 101 2030 102 2034
rect 62 2028 102 2030
rect 62 2024 63 2028
rect 72 2024 74 2028
rect 78 2024 80 2028
rect 84 2024 86 2028
rect 90 2024 92 2028
rect 101 2024 102 2028
rect 62 1768 102 2024
rect 62 1764 63 1768
rect 72 1764 74 1768
rect 78 1764 80 1768
rect 84 1764 86 1768
rect 90 1764 92 1768
rect 101 1764 102 1768
rect 62 1762 102 1764
rect 62 1758 63 1762
rect 72 1758 74 1762
rect 78 1758 80 1762
rect 84 1758 86 1762
rect 90 1758 92 1762
rect 101 1758 102 1762
rect 62 1756 102 1758
rect 62 1752 63 1756
rect 72 1752 74 1756
rect 78 1752 80 1756
rect 84 1752 86 1756
rect 90 1752 92 1756
rect 101 1752 102 1756
rect 62 1750 102 1752
rect 62 1746 63 1750
rect 72 1746 74 1750
rect 78 1746 80 1750
rect 84 1746 86 1750
rect 90 1746 92 1750
rect 101 1746 102 1750
rect 62 1744 102 1746
rect 62 1740 63 1744
rect 72 1740 74 1744
rect 78 1740 80 1744
rect 84 1740 86 1744
rect 90 1740 92 1744
rect 101 1740 102 1744
rect 62 1738 102 1740
rect 62 1734 63 1738
rect 72 1734 74 1738
rect 78 1734 80 1738
rect 84 1734 86 1738
rect 90 1734 92 1738
rect 101 1734 102 1738
rect 62 1732 102 1734
rect 62 1728 63 1732
rect 72 1728 74 1732
rect 78 1728 80 1732
rect 84 1728 86 1732
rect 90 1728 92 1732
rect 101 1728 102 1732
rect 62 1590 102 1728
rect 62 1586 63 1590
rect 72 1586 74 1590
rect 78 1586 80 1590
rect 84 1586 86 1590
rect 90 1586 92 1590
rect 101 1586 102 1590
rect 62 1584 102 1586
rect 62 1580 63 1584
rect 72 1580 74 1584
rect 78 1580 80 1584
rect 84 1580 86 1584
rect 90 1580 92 1584
rect 101 1580 102 1584
rect 62 1578 102 1580
rect 62 1574 63 1578
rect 72 1574 74 1578
rect 78 1574 80 1578
rect 84 1574 86 1578
rect 90 1574 92 1578
rect 101 1574 102 1578
rect 62 1572 102 1574
rect 62 1568 63 1572
rect 72 1568 74 1572
rect 78 1568 80 1572
rect 84 1568 86 1572
rect 90 1568 92 1572
rect 101 1568 102 1572
rect 62 1566 102 1568
rect 62 1562 63 1566
rect 72 1562 74 1566
rect 78 1562 80 1566
rect 84 1562 86 1566
rect 90 1562 92 1566
rect 101 1562 102 1566
rect 62 1560 102 1562
rect 62 1556 63 1560
rect 72 1556 74 1560
rect 78 1556 80 1560
rect 84 1556 86 1560
rect 90 1556 92 1560
rect 101 1556 102 1560
rect 62 1554 102 1556
rect 62 1550 63 1554
rect 72 1550 74 1554
rect 78 1550 80 1554
rect 84 1550 86 1554
rect 90 1550 92 1554
rect 101 1550 102 1554
rect 62 1294 102 1550
rect 62 1290 63 1294
rect 72 1290 74 1294
rect 78 1290 80 1294
rect 84 1290 86 1294
rect 90 1290 92 1294
rect 101 1290 102 1294
rect 62 1288 102 1290
rect 62 1284 63 1288
rect 72 1284 74 1288
rect 78 1284 80 1288
rect 84 1284 86 1288
rect 90 1284 92 1288
rect 101 1284 102 1288
rect 62 1282 102 1284
rect 62 1278 63 1282
rect 72 1278 74 1282
rect 78 1278 80 1282
rect 84 1278 86 1282
rect 90 1278 92 1282
rect 101 1278 102 1282
rect 62 1276 102 1278
rect 62 1272 63 1276
rect 72 1272 74 1276
rect 78 1272 80 1276
rect 84 1272 86 1276
rect 90 1272 92 1276
rect 101 1272 102 1276
rect 62 1270 102 1272
rect 62 1266 63 1270
rect 72 1266 74 1270
rect 78 1266 80 1270
rect 84 1266 86 1270
rect 90 1266 92 1270
rect 101 1266 102 1270
rect 62 1264 102 1266
rect 62 1260 63 1264
rect 72 1260 74 1264
rect 78 1260 80 1264
rect 84 1260 86 1264
rect 90 1260 92 1264
rect 101 1260 102 1264
rect 62 1258 102 1260
rect 62 1254 63 1258
rect 72 1254 74 1258
rect 78 1254 80 1258
rect 84 1254 86 1258
rect 90 1254 92 1258
rect 101 1254 102 1258
rect 62 1116 102 1254
rect 62 1112 63 1116
rect 72 1112 74 1116
rect 78 1112 80 1116
rect 84 1112 86 1116
rect 90 1112 92 1116
rect 101 1112 102 1116
rect 62 1110 102 1112
rect 62 1106 63 1110
rect 72 1106 74 1110
rect 78 1106 80 1110
rect 84 1106 86 1110
rect 90 1106 92 1110
rect 101 1106 102 1110
rect 62 1104 102 1106
rect 62 1100 63 1104
rect 72 1100 74 1104
rect 78 1100 80 1104
rect 84 1100 86 1104
rect 90 1100 92 1104
rect 101 1100 102 1104
rect 62 1098 102 1100
rect 62 1094 63 1098
rect 72 1094 74 1098
rect 78 1094 80 1098
rect 84 1094 86 1098
rect 90 1094 92 1098
rect 101 1094 102 1098
rect 62 1092 102 1094
rect 62 1088 63 1092
rect 72 1088 74 1092
rect 78 1088 80 1092
rect 84 1088 86 1092
rect 90 1088 92 1092
rect 101 1088 102 1092
rect 62 1086 102 1088
rect 62 1082 63 1086
rect 72 1082 74 1086
rect 78 1082 80 1086
rect 84 1082 86 1086
rect 90 1082 92 1086
rect 101 1082 102 1086
rect 62 1080 102 1082
rect 62 1076 63 1080
rect 72 1076 74 1080
rect 78 1076 80 1080
rect 84 1076 86 1080
rect 90 1076 92 1080
rect 101 1076 102 1080
rect 62 820 102 1076
rect 62 816 63 820
rect 72 816 74 820
rect 78 816 80 820
rect 84 816 86 820
rect 90 816 92 820
rect 101 816 102 820
rect 62 814 102 816
rect 62 810 63 814
rect 72 810 74 814
rect 78 810 80 814
rect 84 810 86 814
rect 90 810 92 814
rect 101 810 102 814
rect 62 808 102 810
rect 62 804 63 808
rect 72 804 74 808
rect 78 804 80 808
rect 84 804 86 808
rect 90 804 92 808
rect 101 804 102 808
rect 62 802 102 804
rect 62 798 63 802
rect 72 798 74 802
rect 78 798 80 802
rect 84 798 86 802
rect 90 798 92 802
rect 101 798 102 802
rect 62 796 102 798
rect 62 792 63 796
rect 72 792 74 796
rect 78 792 80 796
rect 84 792 86 796
rect 90 792 92 796
rect 101 792 102 796
rect 62 790 102 792
rect 62 786 63 790
rect 72 786 74 790
rect 78 786 80 790
rect 84 786 86 790
rect 90 786 92 790
rect 101 786 102 790
rect 62 784 102 786
rect 62 780 63 784
rect 72 780 74 784
rect 78 780 80 784
rect 84 780 86 784
rect 90 780 92 784
rect 101 780 102 784
rect 62 642 102 780
rect 62 638 63 642
rect 72 638 74 642
rect 78 638 80 642
rect 84 638 86 642
rect 90 638 92 642
rect 101 638 102 642
rect 62 636 102 638
rect 62 632 63 636
rect 72 632 74 636
rect 78 632 80 636
rect 84 632 86 636
rect 90 632 92 636
rect 101 632 102 636
rect 62 630 102 632
rect 62 626 63 630
rect 72 626 74 630
rect 78 626 80 630
rect 84 626 86 630
rect 90 626 92 630
rect 101 626 102 630
rect 62 624 102 626
rect 62 620 63 624
rect 72 620 74 624
rect 78 620 80 624
rect 84 620 86 624
rect 90 620 92 624
rect 101 620 102 624
rect 62 618 102 620
rect 62 614 63 618
rect 72 614 74 618
rect 78 614 80 618
rect 84 614 86 618
rect 90 614 92 618
rect 101 614 102 618
rect 62 612 102 614
rect 62 608 63 612
rect 72 608 74 612
rect 78 608 80 612
rect 84 608 86 612
rect 90 608 92 612
rect 101 608 102 612
rect 62 606 102 608
rect 62 602 63 606
rect 72 602 74 606
rect 78 602 80 606
rect 84 602 86 606
rect 90 602 92 606
rect 101 602 102 606
rect 62 346 102 602
rect 62 342 63 346
rect 72 342 74 346
rect 78 342 80 346
rect 84 342 86 346
rect 90 342 92 346
rect 101 342 102 346
rect 62 340 102 342
rect 62 336 63 340
rect 72 336 74 340
rect 78 336 80 340
rect 84 336 86 340
rect 90 336 92 340
rect 101 336 102 340
rect 62 334 102 336
rect 62 330 63 334
rect 72 330 74 334
rect 78 330 80 334
rect 84 330 86 334
rect 90 330 92 334
rect 101 330 102 334
rect 62 328 102 330
rect 62 324 63 328
rect 72 324 74 328
rect 78 324 80 328
rect 84 324 86 328
rect 90 324 92 328
rect 101 324 102 328
rect 62 322 102 324
rect 62 318 63 322
rect 72 318 74 322
rect 78 318 80 322
rect 84 318 86 322
rect 90 318 92 322
rect 101 318 102 322
rect 62 316 102 318
rect 62 312 63 316
rect 72 312 74 316
rect 78 312 80 316
rect 84 312 86 316
rect 90 312 92 316
rect 101 312 102 316
rect 62 310 102 312
rect 62 306 63 310
rect 72 306 74 310
rect 78 306 80 310
rect 84 306 86 310
rect 90 306 92 310
rect 101 306 102 310
rect 62 168 102 306
rect 62 164 63 168
rect 72 164 74 168
rect 78 164 80 168
rect 84 164 86 168
rect 90 164 92 168
rect 101 164 102 168
rect 62 162 102 164
rect 62 158 63 162
rect 72 158 74 162
rect 78 158 80 162
rect 84 158 86 162
rect 90 158 92 162
rect 101 158 102 162
rect 62 156 102 158
rect 62 152 63 156
rect 72 152 74 156
rect 78 152 80 156
rect 84 152 86 156
rect 90 152 92 156
rect 101 152 102 156
rect 62 150 102 152
rect 62 146 63 150
rect 72 146 74 150
rect 78 146 80 150
rect 84 146 86 150
rect 90 146 92 150
rect 101 146 102 150
rect 62 144 102 146
rect 62 140 63 144
rect 72 140 74 144
rect 78 140 80 144
rect 84 140 86 144
rect 90 140 92 144
rect 101 140 102 144
rect 62 138 102 140
rect 62 134 63 138
rect 72 134 74 138
rect 78 134 80 138
rect 84 134 86 138
rect 90 134 92 138
rect 101 134 102 138
rect 62 132 102 134
rect 62 128 63 132
rect 72 128 74 132
rect 78 128 80 132
rect 84 128 86 132
rect 90 128 92 132
rect 101 128 102 132
rect 62 84 102 128
rect 106 4094 146 4226
rect 106 4090 107 4094
rect 111 4090 119 4094
rect 123 4090 146 4094
rect 106 4088 146 4090
rect 106 4084 107 4088
rect 111 4084 119 4088
rect 123 4084 131 4088
rect 135 4084 146 4088
rect 106 4082 146 4084
rect 106 4078 107 4082
rect 111 4078 119 4082
rect 123 4078 131 4082
rect 135 4078 146 4082
rect 106 4076 146 4078
rect 106 4072 107 4076
rect 111 4072 119 4076
rect 123 4072 131 4076
rect 135 4072 146 4076
rect 106 4070 146 4072
rect 106 4066 107 4070
rect 111 4066 119 4070
rect 123 4066 131 4070
rect 135 4066 146 4070
rect 106 4064 146 4066
rect 106 4060 107 4064
rect 111 4060 119 4064
rect 123 4060 131 4064
rect 135 4060 146 4064
rect 106 4058 146 4060
rect 106 4054 107 4058
rect 111 4054 119 4058
rect 123 4054 131 4058
rect 135 4054 146 4058
rect 106 4004 146 4054
rect 106 4000 107 4004
rect 111 4000 119 4004
rect 123 4000 131 4004
rect 135 4000 146 4004
rect 106 3998 146 4000
rect 106 3994 107 3998
rect 111 3994 119 3998
rect 123 3994 131 3998
rect 135 3994 146 3998
rect 106 3992 146 3994
rect 106 3988 107 3992
rect 111 3988 119 3992
rect 123 3988 131 3992
rect 135 3988 146 3992
rect 106 3986 146 3988
rect 106 3982 107 3986
rect 111 3982 119 3986
rect 123 3982 131 3986
rect 135 3982 146 3986
rect 106 3980 146 3982
rect 106 3976 107 3980
rect 111 3976 119 3980
rect 123 3976 131 3980
rect 135 3976 146 3980
rect 106 3974 146 3976
rect 106 3970 107 3974
rect 111 3970 119 3974
rect 123 3970 131 3974
rect 135 3970 146 3974
rect 106 3968 146 3970
rect 106 3964 107 3968
rect 111 3964 119 3968
rect 123 3964 146 3968
rect 106 3620 146 3964
rect 106 3616 107 3620
rect 111 3616 119 3620
rect 123 3616 146 3620
rect 106 3614 146 3616
rect 106 3610 107 3614
rect 111 3610 119 3614
rect 123 3610 131 3614
rect 135 3610 146 3614
rect 106 3608 146 3610
rect 106 3604 107 3608
rect 111 3604 119 3608
rect 123 3604 131 3608
rect 135 3604 146 3608
rect 106 3602 146 3604
rect 106 3598 107 3602
rect 111 3598 119 3602
rect 123 3598 131 3602
rect 135 3598 146 3602
rect 106 3596 146 3598
rect 106 3592 107 3596
rect 111 3592 119 3596
rect 123 3592 131 3596
rect 135 3592 146 3596
rect 106 3590 146 3592
rect 106 3586 107 3590
rect 111 3586 119 3590
rect 123 3586 131 3590
rect 135 3586 146 3590
rect 106 3584 146 3586
rect 106 3580 107 3584
rect 111 3580 119 3584
rect 123 3580 131 3584
rect 135 3580 146 3584
rect 106 3530 146 3580
rect 106 3526 107 3530
rect 111 3526 119 3530
rect 123 3526 131 3530
rect 135 3526 146 3530
rect 106 3524 146 3526
rect 106 3520 107 3524
rect 111 3520 119 3524
rect 123 3520 131 3524
rect 135 3520 146 3524
rect 106 3518 146 3520
rect 106 3514 107 3518
rect 111 3514 119 3518
rect 123 3514 131 3518
rect 135 3514 146 3518
rect 106 3512 146 3514
rect 106 3508 107 3512
rect 111 3508 119 3512
rect 123 3508 131 3512
rect 135 3508 146 3512
rect 106 3506 146 3508
rect 106 3502 107 3506
rect 111 3502 119 3506
rect 123 3502 131 3506
rect 135 3502 146 3506
rect 106 3500 146 3502
rect 106 3496 107 3500
rect 111 3496 119 3500
rect 123 3496 131 3500
rect 135 3496 146 3500
rect 106 3494 146 3496
rect 106 3490 107 3494
rect 111 3490 119 3494
rect 123 3490 146 3494
rect 106 3146 146 3490
rect 106 3142 107 3146
rect 111 3142 119 3146
rect 123 3142 146 3146
rect 106 3140 146 3142
rect 106 3136 107 3140
rect 111 3136 119 3140
rect 123 3136 131 3140
rect 135 3136 146 3140
rect 106 3134 146 3136
rect 106 3130 107 3134
rect 111 3130 119 3134
rect 123 3130 131 3134
rect 135 3130 146 3134
rect 106 3128 146 3130
rect 106 3124 107 3128
rect 111 3124 119 3128
rect 123 3124 131 3128
rect 135 3124 146 3128
rect 106 3122 146 3124
rect 106 3118 107 3122
rect 111 3118 119 3122
rect 123 3118 131 3122
rect 135 3118 146 3122
rect 106 3116 146 3118
rect 106 3112 107 3116
rect 111 3112 119 3116
rect 123 3112 131 3116
rect 135 3112 146 3116
rect 106 3110 146 3112
rect 106 3106 107 3110
rect 111 3106 119 3110
rect 123 3106 131 3110
rect 135 3106 146 3110
rect 106 3056 146 3106
rect 106 3052 107 3056
rect 111 3052 119 3056
rect 123 3052 131 3056
rect 135 3052 146 3056
rect 106 3050 146 3052
rect 106 3046 107 3050
rect 111 3046 119 3050
rect 123 3046 131 3050
rect 135 3046 146 3050
rect 106 3044 146 3046
rect 106 3040 107 3044
rect 111 3040 119 3044
rect 123 3040 131 3044
rect 135 3040 146 3044
rect 106 3038 146 3040
rect 106 3034 107 3038
rect 111 3034 119 3038
rect 123 3034 131 3038
rect 135 3034 146 3038
rect 106 3032 146 3034
rect 106 3028 107 3032
rect 111 3028 119 3032
rect 123 3028 131 3032
rect 135 3028 146 3032
rect 106 3026 146 3028
rect 106 3022 107 3026
rect 111 3022 119 3026
rect 123 3022 131 3026
rect 135 3022 146 3026
rect 106 3020 146 3022
rect 106 3016 107 3020
rect 111 3016 119 3020
rect 123 3016 146 3020
rect 106 2672 146 3016
rect 106 2668 107 2672
rect 111 2668 119 2672
rect 123 2668 146 2672
rect 106 2666 146 2668
rect 106 2662 107 2666
rect 111 2662 119 2666
rect 123 2662 131 2666
rect 135 2662 146 2666
rect 106 2660 146 2662
rect 106 2656 107 2660
rect 111 2656 119 2660
rect 123 2656 131 2660
rect 135 2656 146 2660
rect 106 2654 146 2656
rect 106 2650 107 2654
rect 111 2650 119 2654
rect 123 2650 131 2654
rect 135 2650 146 2654
rect 106 2648 146 2650
rect 106 2644 107 2648
rect 111 2644 119 2648
rect 123 2644 131 2648
rect 135 2644 146 2648
rect 106 2642 146 2644
rect 106 2638 107 2642
rect 111 2638 119 2642
rect 123 2638 131 2642
rect 135 2638 146 2642
rect 106 2636 146 2638
rect 106 2632 107 2636
rect 111 2632 119 2636
rect 123 2632 131 2636
rect 135 2632 146 2636
rect 106 2582 146 2632
rect 106 2578 107 2582
rect 111 2578 119 2582
rect 123 2578 131 2582
rect 135 2578 146 2582
rect 106 2576 146 2578
rect 106 2572 107 2576
rect 111 2572 119 2576
rect 123 2572 131 2576
rect 135 2572 146 2576
rect 106 2570 146 2572
rect 106 2566 107 2570
rect 111 2566 119 2570
rect 123 2566 131 2570
rect 135 2566 146 2570
rect 106 2564 146 2566
rect 106 2560 107 2564
rect 111 2560 119 2564
rect 123 2560 131 2564
rect 135 2560 146 2564
rect 106 2558 146 2560
rect 106 2554 107 2558
rect 111 2554 119 2558
rect 123 2554 131 2558
rect 135 2554 146 2558
rect 106 2552 146 2554
rect 106 2548 107 2552
rect 111 2548 119 2552
rect 123 2548 131 2552
rect 135 2548 146 2552
rect 106 2546 146 2548
rect 106 2542 107 2546
rect 111 2542 119 2546
rect 123 2542 146 2546
rect 106 2198 146 2542
rect 106 2194 107 2198
rect 111 2194 119 2198
rect 123 2194 146 2198
rect 106 2192 146 2194
rect 106 2188 107 2192
rect 111 2188 119 2192
rect 123 2188 131 2192
rect 135 2188 146 2192
rect 106 2186 146 2188
rect 106 2182 107 2186
rect 111 2182 119 2186
rect 123 2182 131 2186
rect 135 2182 146 2186
rect 106 2180 146 2182
rect 106 2176 107 2180
rect 111 2176 119 2180
rect 123 2176 131 2180
rect 135 2176 146 2180
rect 106 2174 146 2176
rect 106 2170 107 2174
rect 111 2170 119 2174
rect 123 2170 131 2174
rect 135 2170 146 2174
rect 106 2168 146 2170
rect 106 2164 107 2168
rect 111 2164 119 2168
rect 123 2164 131 2168
rect 135 2164 146 2168
rect 106 2162 146 2164
rect 106 2158 107 2162
rect 111 2158 119 2162
rect 123 2158 131 2162
rect 135 2158 146 2162
rect 106 2108 146 2158
rect 106 2104 107 2108
rect 111 2104 119 2108
rect 123 2104 131 2108
rect 135 2104 146 2108
rect 106 2102 146 2104
rect 106 2098 107 2102
rect 111 2098 119 2102
rect 123 2098 131 2102
rect 135 2098 146 2102
rect 106 2096 146 2098
rect 106 2092 107 2096
rect 111 2092 119 2096
rect 123 2092 131 2096
rect 135 2092 146 2096
rect 106 2090 146 2092
rect 106 2086 107 2090
rect 111 2086 119 2090
rect 123 2086 131 2090
rect 135 2086 146 2090
rect 106 2084 146 2086
rect 106 2080 107 2084
rect 111 2080 119 2084
rect 123 2080 131 2084
rect 135 2080 146 2084
rect 106 2078 146 2080
rect 106 2074 107 2078
rect 111 2074 119 2078
rect 123 2074 131 2078
rect 135 2074 146 2078
rect 106 2072 146 2074
rect 106 2068 107 2072
rect 111 2068 119 2072
rect 123 2068 146 2072
rect 106 1724 146 2068
rect 106 1720 107 1724
rect 111 1720 119 1724
rect 123 1720 146 1724
rect 106 1718 146 1720
rect 106 1714 107 1718
rect 111 1714 119 1718
rect 123 1714 131 1718
rect 135 1714 146 1718
rect 106 1712 146 1714
rect 106 1708 107 1712
rect 111 1708 119 1712
rect 123 1708 131 1712
rect 135 1708 146 1712
rect 106 1706 146 1708
rect 106 1702 107 1706
rect 111 1702 119 1706
rect 123 1702 131 1706
rect 135 1702 146 1706
rect 106 1700 146 1702
rect 106 1696 107 1700
rect 111 1696 119 1700
rect 123 1696 131 1700
rect 135 1696 146 1700
rect 106 1694 146 1696
rect 106 1690 107 1694
rect 111 1690 119 1694
rect 123 1690 131 1694
rect 135 1690 146 1694
rect 106 1688 146 1690
rect 106 1684 107 1688
rect 111 1684 119 1688
rect 123 1684 131 1688
rect 135 1684 146 1688
rect 106 1634 146 1684
rect 106 1630 107 1634
rect 111 1630 119 1634
rect 123 1630 131 1634
rect 135 1630 146 1634
rect 106 1628 146 1630
rect 106 1624 107 1628
rect 111 1624 119 1628
rect 123 1624 131 1628
rect 135 1624 146 1628
rect 106 1622 146 1624
rect 106 1618 107 1622
rect 111 1618 119 1622
rect 123 1618 131 1622
rect 135 1618 146 1622
rect 106 1616 146 1618
rect 106 1612 107 1616
rect 111 1612 119 1616
rect 123 1612 131 1616
rect 135 1612 146 1616
rect 106 1610 146 1612
rect 106 1606 107 1610
rect 111 1606 119 1610
rect 123 1606 131 1610
rect 135 1606 146 1610
rect 106 1604 146 1606
rect 106 1600 107 1604
rect 111 1600 119 1604
rect 123 1600 131 1604
rect 135 1600 146 1604
rect 106 1598 146 1600
rect 106 1594 107 1598
rect 111 1594 119 1598
rect 123 1594 146 1598
rect 106 1250 146 1594
rect 106 1246 107 1250
rect 111 1246 119 1250
rect 123 1246 146 1250
rect 106 1244 146 1246
rect 106 1240 107 1244
rect 111 1240 119 1244
rect 123 1240 131 1244
rect 135 1240 146 1244
rect 106 1238 146 1240
rect 106 1234 107 1238
rect 111 1234 119 1238
rect 123 1234 131 1238
rect 135 1234 146 1238
rect 106 1232 146 1234
rect 106 1228 107 1232
rect 111 1228 119 1232
rect 123 1228 131 1232
rect 135 1228 146 1232
rect 106 1226 146 1228
rect 106 1222 107 1226
rect 111 1222 119 1226
rect 123 1222 131 1226
rect 135 1222 146 1226
rect 106 1220 146 1222
rect 106 1216 107 1220
rect 111 1216 119 1220
rect 123 1216 131 1220
rect 135 1216 146 1220
rect 106 1214 146 1216
rect 106 1210 107 1214
rect 111 1210 119 1214
rect 123 1210 131 1214
rect 135 1210 146 1214
rect 106 1160 146 1210
rect 106 1156 107 1160
rect 111 1156 119 1160
rect 123 1156 131 1160
rect 135 1156 146 1160
rect 106 1154 146 1156
rect 106 1150 107 1154
rect 111 1150 119 1154
rect 123 1150 131 1154
rect 135 1150 146 1154
rect 106 1148 146 1150
rect 106 1144 107 1148
rect 111 1144 119 1148
rect 123 1144 131 1148
rect 135 1144 146 1148
rect 106 1142 146 1144
rect 106 1138 107 1142
rect 111 1138 119 1142
rect 123 1138 131 1142
rect 135 1138 146 1142
rect 106 1136 146 1138
rect 106 1132 107 1136
rect 111 1132 119 1136
rect 123 1132 131 1136
rect 135 1132 146 1136
rect 106 1130 146 1132
rect 106 1126 107 1130
rect 111 1126 119 1130
rect 123 1126 131 1130
rect 135 1126 146 1130
rect 106 1124 146 1126
rect 106 1120 107 1124
rect 111 1120 119 1124
rect 123 1120 146 1124
rect 106 776 146 1120
rect 106 772 107 776
rect 111 772 119 776
rect 123 772 146 776
rect 106 770 146 772
rect 106 766 107 770
rect 111 766 119 770
rect 123 766 131 770
rect 135 766 146 770
rect 106 764 146 766
rect 106 760 107 764
rect 111 760 119 764
rect 123 760 131 764
rect 135 760 146 764
rect 106 758 146 760
rect 106 754 107 758
rect 111 754 119 758
rect 123 754 131 758
rect 135 754 146 758
rect 106 752 146 754
rect 106 748 107 752
rect 111 748 119 752
rect 123 748 131 752
rect 135 748 146 752
rect 106 746 146 748
rect 106 742 107 746
rect 111 742 119 746
rect 123 742 131 746
rect 135 742 146 746
rect 106 740 146 742
rect 106 736 107 740
rect 111 736 119 740
rect 123 736 131 740
rect 135 736 146 740
rect 106 686 146 736
rect 106 682 107 686
rect 111 682 119 686
rect 123 682 131 686
rect 135 682 146 686
rect 106 680 146 682
rect 106 676 107 680
rect 111 676 119 680
rect 123 676 131 680
rect 135 676 146 680
rect 106 674 146 676
rect 106 670 107 674
rect 111 670 119 674
rect 123 670 131 674
rect 135 670 146 674
rect 106 668 146 670
rect 106 664 107 668
rect 111 664 119 668
rect 123 664 131 668
rect 135 664 146 668
rect 106 662 146 664
rect 106 658 107 662
rect 111 658 119 662
rect 123 658 131 662
rect 135 658 146 662
rect 106 656 146 658
rect 106 652 107 656
rect 111 652 119 656
rect 123 652 131 656
rect 135 652 146 656
rect 106 650 146 652
rect 106 646 107 650
rect 111 646 119 650
rect 123 646 146 650
rect 106 302 146 646
rect 106 298 107 302
rect 111 298 119 302
rect 123 298 146 302
rect 106 296 146 298
rect 106 292 107 296
rect 111 292 119 296
rect 123 292 131 296
rect 135 292 146 296
rect 106 290 146 292
rect 106 286 107 290
rect 111 286 119 290
rect 123 286 131 290
rect 135 286 146 290
rect 106 284 146 286
rect 106 280 107 284
rect 111 280 119 284
rect 123 280 131 284
rect 135 280 146 284
rect 106 278 146 280
rect 106 274 107 278
rect 111 274 119 278
rect 123 274 131 278
rect 135 274 146 278
rect 106 272 146 274
rect 106 268 107 272
rect 111 268 119 272
rect 123 268 131 272
rect 135 268 146 272
rect 106 266 146 268
rect 106 262 107 266
rect 111 262 119 266
rect 123 262 131 266
rect 135 262 146 266
rect 106 212 146 262
rect 106 208 107 212
rect 111 208 119 212
rect 123 208 131 212
rect 135 208 146 212
rect 106 206 146 208
rect 106 202 107 206
rect 111 202 119 206
rect 123 202 131 206
rect 135 202 146 206
rect 106 200 146 202
rect 106 196 107 200
rect 111 196 119 200
rect 123 196 131 200
rect 135 196 146 200
rect 106 194 146 196
rect 106 190 107 194
rect 111 190 119 194
rect 123 190 131 194
rect 135 190 146 194
rect 106 188 146 190
rect 106 184 107 188
rect 111 184 119 188
rect 123 184 131 188
rect 135 184 146 188
rect 106 182 146 184
rect 106 178 107 182
rect 111 178 119 182
rect 123 178 131 182
rect 135 178 146 182
rect 106 176 146 178
rect 106 172 107 176
rect 111 172 119 176
rect 123 172 146 176
rect 106 117 146 172
rect 106 113 107 117
rect 111 113 113 117
rect 117 113 119 117
rect 123 113 125 117
rect 129 113 131 117
rect 135 113 146 117
rect 106 111 146 113
rect 106 107 107 111
rect 111 107 113 111
rect 117 107 119 111
rect 123 107 125 111
rect 129 107 131 111
rect 135 107 146 111
rect 106 105 146 107
rect 106 101 107 105
rect 111 101 113 105
rect 117 101 119 105
rect 123 101 125 105
rect 129 101 131 105
rect 135 101 146 105
rect 106 99 146 101
rect 106 95 107 99
rect 111 95 113 99
rect 117 95 119 99
rect 123 95 125 99
rect 129 95 131 99
rect 135 95 146 99
rect 106 93 146 95
rect 106 89 107 93
rect 111 89 113 93
rect 117 89 119 93
rect 123 89 125 93
rect 129 89 131 93
rect 135 89 146 93
rect 106 87 146 89
rect 106 83 107 87
rect 111 83 113 87
rect 117 83 119 87
rect 123 83 125 87
rect 129 83 131 87
rect 135 83 146 87
rect 106 81 146 83
rect 106 77 107 81
rect 111 77 113 81
rect 117 77 119 81
rect 123 77 125 81
rect 129 77 131 81
rect 135 77 146 81
rect 106 75 146 77
rect 106 71 107 75
rect 111 71 113 75
rect 117 71 119 75
rect 123 71 125 75
rect 129 71 131 75
rect 135 71 146 75
rect 106 69 146 71
rect 106 65 107 69
rect 111 65 113 69
rect 117 65 119 69
rect 123 65 125 69
rect 129 65 131 69
rect 135 65 146 69
rect 106 63 146 65
rect 106 59 107 63
rect 111 59 113 63
rect 117 59 119 63
rect 123 59 125 63
rect 129 59 131 63
rect 135 59 146 63
rect 106 57 146 59
rect 106 53 107 57
rect 111 53 113 57
rect 117 53 119 57
rect 123 53 125 57
rect 129 53 131 57
rect 135 53 146 57
rect 106 51 146 53
rect 106 47 107 51
rect 111 47 113 51
rect 117 47 119 51
rect 123 47 125 51
rect 129 47 131 51
rect 135 47 146 51
rect 106 40 146 47
<< m3contact >>
rect 107 113 111 117
rect 113 113 117 117
rect 119 113 123 117
rect 125 113 129 117
rect 131 113 135 117
rect 107 107 111 111
rect 113 107 117 111
rect 119 107 123 111
rect 125 107 129 111
rect 131 107 135 111
rect 107 101 111 105
rect 113 101 117 105
rect 119 101 123 105
rect 125 101 129 105
rect 131 101 135 105
rect 107 95 111 99
rect 113 95 117 99
rect 119 95 123 99
rect 125 95 129 99
rect 131 95 135 99
rect 107 89 111 93
rect 113 89 117 93
rect 119 89 123 93
rect 125 89 129 93
rect 131 89 135 93
rect 107 83 111 87
rect 113 83 117 87
rect 119 83 123 87
rect 125 83 129 87
rect 131 83 135 87
rect 107 77 111 81
rect 113 77 117 81
rect 119 77 123 81
rect 125 77 129 81
rect 131 77 135 81
rect 107 71 111 75
rect 113 71 117 75
rect 119 71 123 75
rect 125 71 129 75
rect 131 71 135 75
rect 107 65 111 69
rect 113 65 117 69
rect 119 65 123 69
rect 125 65 129 69
rect 131 65 135 69
rect 107 59 111 63
rect 113 59 117 63
rect 119 59 123 63
rect 125 59 129 63
rect 131 59 135 63
rect 107 53 111 57
rect 113 53 117 57
rect 119 53 123 57
rect 125 53 129 57
rect 131 53 135 57
rect 107 47 111 51
rect 113 47 117 51
rect 119 47 123 51
rect 125 47 129 51
rect 131 47 135 51
<< metal3 >>
rect 106 117 137 118
rect 106 113 107 117
rect 111 113 113 117
rect 117 113 119 117
rect 123 113 125 117
rect 129 113 131 117
rect 135 113 137 117
rect 106 111 137 113
rect 106 107 107 111
rect 111 107 113 111
rect 117 107 119 111
rect 123 107 125 111
rect 129 107 131 111
rect 135 107 137 111
rect 106 105 137 107
rect 106 101 107 105
rect 111 101 113 105
rect 117 101 119 105
rect 123 101 125 105
rect 129 101 131 105
rect 135 101 137 105
rect 106 99 137 101
rect 106 95 107 99
rect 111 95 113 99
rect 117 95 119 99
rect 123 95 125 99
rect 129 95 131 99
rect 135 95 137 99
rect 106 93 137 95
rect 106 89 107 93
rect 111 89 113 93
rect 117 89 119 93
rect 123 89 125 93
rect 129 89 131 93
rect 135 89 137 93
rect 106 87 137 89
rect 106 83 107 87
rect 111 83 113 87
rect 117 83 119 87
rect 123 83 125 87
rect 129 83 131 87
rect 135 83 137 87
rect 106 81 137 83
rect 106 77 107 81
rect 111 77 113 81
rect 117 77 119 81
rect 123 77 125 81
rect 129 77 131 81
rect 135 77 137 81
rect 106 75 137 77
rect 106 71 107 75
rect 111 71 113 75
rect 117 71 119 75
rect 123 71 125 75
rect 129 71 131 75
rect 135 71 137 75
rect 106 69 137 71
rect 106 65 107 69
rect 111 65 113 69
rect 117 65 119 69
rect 123 65 125 69
rect 129 65 131 69
rect 135 65 137 69
rect 106 63 137 65
rect 106 59 107 63
rect 111 59 113 63
rect 117 59 119 63
rect 123 59 125 63
rect 129 59 131 63
rect 135 59 137 63
rect 106 57 137 59
rect 106 53 107 57
rect 111 53 113 57
rect 117 53 119 57
rect 123 53 125 57
rect 129 53 131 57
rect 135 53 137 57
rect 106 51 137 53
rect 106 47 107 51
rect 111 47 113 51
rect 117 47 119 51
rect 123 47 125 51
rect 129 47 131 51
rect 135 47 137 51
rect 106 40 137 47
<< labels >>
rlabel m2contact 0 326 0 326 4 Gnd
rlabel m2contact 0 192 0 192 4 CVdd
rlabel m2contact 0 220 0 220 4 Bias
rlabel m2contact 0 253 0 253 4 Bias
rlabel m2contact 0 282 0 282 4 CVdd
rlabel m2contact 0 800 0 800 4 Gnd
rlabel m2contact 0 622 0 622 4 Gnd
rlabel m2contact 0 666 0 666 4 CVdd
rlabel m2contact 0 694 0 694 4 Bias
rlabel m2contact 0 727 0 727 4 Bias
rlabel m2contact 0 756 0 756 4 CVdd
rlabel m2contact 0 1274 0 1274 4 Gnd
rlabel m2contact 0 1096 0 1096 4 Gnd
rlabel m2contact 0 1140 0 1140 4 CVdd
rlabel m2contact 0 1168 0 1168 4 Bias
rlabel m2contact 0 1201 0 1201 4 Bias
rlabel m2contact 0 1230 0 1230 4 CVdd
rlabel m2contact 0 1748 0 1748 4 Gnd
rlabel m2contact 0 1570 0 1570 4 Gnd
rlabel m2contact 0 1614 0 1614 4 CVdd
rlabel m2contact 0 1642 0 1642 4 Bias
rlabel m2contact 0 1675 0 1675 4 Bias
rlabel m2contact 0 1704 0 1704 4 CVdd
rlabel m2contact 0 2222 0 2222 4 Gnd
rlabel m2contact 0 2044 0 2044 4 Gnd
rlabel m2contact 0 2088 0 2088 4 CVdd
rlabel m2contact 0 2116 0 2116 4 Bias
rlabel m2contact 0 2149 0 2149 4 Bias
rlabel m2contact 0 2178 0 2178 4 CVdd
rlabel m2contact 0 2696 0 2696 4 Gnd
rlabel m2contact 0 2518 0 2518 4 Gnd
rlabel m2contact 0 2562 0 2562 4 CVdd
rlabel m2contact 0 2590 0 2590 4 Bias
rlabel m2contact 0 2623 0 2623 4 Bias
rlabel m2contact 0 2652 0 2652 4 CVdd
rlabel m2contact 0 3170 0 3170 4 Gnd
rlabel m2contact 0 2992 0 2992 4 Gnd
rlabel m2contact 0 3036 0 3036 4 CVdd
rlabel m2contact 0 3064 0 3064 4 Bias
rlabel m2contact 0 3097 0 3097 4 Bias
rlabel m2contact 0 3126 0 3126 4 CVdd
rlabel m2contact 0 3644 0 3644 4 Gnd
rlabel m2contact 0 3466 0 3466 4 Gnd
rlabel m2contact 0 3510 0 3510 4 CVdd
rlabel m2contact 0 3538 0 3538 4 Bias
rlabel m2contact 0 3571 0 3571 4 Bias
rlabel m2contact 0 3600 0 3600 4 CVdd
rlabel m2contact 0 3940 0 3940 4 Gnd
rlabel m2contact 0 3984 0 3984 4 CVdd
rlabel m2contact 0 4012 0 4012 4 Bias
rlabel m2contact 0 4045 0 4045 4 Bias
rlabel m2contact 0 4074 0 4074 4 CVdd
<< end >>
