magic
tech scmos
timestamp 1413439199
<< nwell >>
rect -6 128 0 130
rect -130 124 11 128
rect -137 120 -133 124
rect -6 97 0 124
rect -6 93 4 97
rect -6 48 0 93
rect 254 82 258 121
<< pwell >>
rect -6 36 2 48
rect -11 17 4 36
rect -6 11 4 17
rect -6 0 2 11
rect -164 -32 -141 -28
rect -144 -38 -22 -34
<< polycontact >>
rect -137 120 -133 124
rect 0 93 4 97
rect -11 32 -7 36
rect 0 32 4 36
rect 0 17 4 21
<< metal1 >>
rect -130 124 11 128
rect -7 93 0 97
rect -11 21 -7 32
rect -11 17 0 21
rect 7 3 127 7
rect -145 -34 -140 -12
rect -7 -25 0 -21
rect 7 -34 11 3
rect -145 -38 11 -34
<< m2contact >>
rect -137 124 -133 128
rect 254 82 258 86
rect 0 28 4 32
rect 0 -25 4 -21
<< metal2 >>
rect -133 124 258 128
rect 254 86 258 124
rect 0 -21 4 28
use bias  bias_0
timestamp 1413439122
transform 1 0 -198 0 1 -29
box -67 -9 192 162
use amp  amp_0
timestamp 1413433214
transform 1 0 7 0 1 72
box -7 -72 252 58
<< end >>
