magic
tech scmos
timestamp 1259953556
<< nwell >>
rect 111 323 155 361
rect 167 323 211 361
rect 311 341 468 361
rect 243 311 468 341
rect 418 159 468 311
<< ntransistor >>
rect 255 347 257 356
rect 260 347 262 356
rect 268 347 270 356
rect 273 347 275 356
rect 281 347 283 356
rect 289 347 291 356
rect 297 347 299 356
rect 424 138 462 140
rect 424 130 462 132
rect 424 122 462 124
rect 424 114 462 116
rect 424 106 462 108
rect 424 98 462 100
rect 424 90 462 92
rect 424 82 462 84
rect 424 74 462 76
rect 424 66 462 68
rect 424 58 462 60
rect 424 50 462 52
rect 424 42 462 44
rect 424 34 462 36
rect 424 26 462 28
rect 424 18 462 20
<< ptransistor >>
rect 255 317 257 335
rect 260 317 262 335
rect 268 317 270 335
rect 273 317 275 335
rect 281 317 283 335
rect 289 317 291 335
rect 297 317 299 335
rect 326 317 328 355
rect 334 317 336 355
rect 342 317 344 355
rect 350 317 352 355
rect 358 317 360 355
rect 366 317 368 355
rect 374 317 376 355
rect 382 317 384 355
rect 390 317 392 355
rect 398 317 400 355
rect 406 317 408 355
rect 414 317 416 355
rect 422 317 424 355
rect 430 317 432 355
rect 438 317 440 355
rect 446 317 448 355
rect 424 294 462 296
rect 424 286 462 288
rect 424 278 462 280
rect 424 270 462 272
rect 424 262 462 264
rect 424 254 462 256
rect 424 246 462 248
rect 424 238 462 240
rect 424 230 462 232
rect 424 222 462 224
rect 424 214 462 216
rect 424 206 462 208
rect 424 198 462 200
rect 424 190 462 192
rect 424 182 462 184
rect 424 174 462 176
<< ndiffusion >>
rect 34 359 46 360
rect 34 355 35 359
rect 39 355 41 359
rect 45 355 46 359
rect 34 353 46 355
rect 34 349 35 353
rect 39 349 41 353
rect 45 349 46 353
rect 34 347 46 349
rect 34 343 35 347
rect 39 343 41 347
rect 45 343 46 347
rect 34 341 46 343
rect 34 337 35 341
rect 39 337 41 341
rect 45 337 46 341
rect 34 335 46 337
rect 34 331 35 335
rect 39 331 41 335
rect 45 331 46 335
rect 34 329 46 331
rect 34 325 35 329
rect 39 325 41 329
rect 45 325 46 329
rect 34 324 46 325
rect 60 359 72 360
rect 60 355 61 359
rect 65 355 67 359
rect 71 355 72 359
rect 60 353 72 355
rect 60 349 61 353
rect 65 349 67 353
rect 71 349 72 353
rect 60 347 72 349
rect 60 343 61 347
rect 65 343 67 347
rect 71 343 72 347
rect 60 341 72 343
rect 60 337 61 341
rect 65 337 67 341
rect 71 337 72 341
rect 60 335 72 337
rect 60 331 61 335
rect 65 331 67 335
rect 71 331 72 335
rect 60 329 72 331
rect 60 325 61 329
rect 65 325 67 329
rect 71 325 72 329
rect 60 324 72 325
rect 86 359 98 360
rect 86 355 87 359
rect 91 355 93 359
rect 97 355 98 359
rect 86 353 98 355
rect 86 349 87 353
rect 91 349 93 353
rect 97 349 98 353
rect 86 347 98 349
rect 86 343 87 347
rect 91 343 93 347
rect 97 343 98 347
rect 86 341 98 343
rect 86 337 87 341
rect 91 337 93 341
rect 97 337 98 341
rect 86 335 98 337
rect 86 331 87 335
rect 91 331 93 335
rect 97 331 98 335
rect 86 329 98 331
rect 86 325 87 329
rect 91 325 93 329
rect 97 325 98 329
rect 86 324 98 325
rect 249 355 255 356
rect 249 351 250 355
rect 254 351 255 355
rect 249 347 255 351
rect 257 347 260 356
rect 262 352 268 356
rect 262 348 263 352
rect 267 348 268 352
rect 262 347 268 348
rect 270 347 273 356
rect 275 355 281 356
rect 275 351 276 355
rect 280 351 281 355
rect 275 347 281 351
rect 283 352 289 356
rect 283 348 284 352
rect 288 348 289 352
rect 283 347 289 348
rect 291 355 297 356
rect 291 351 292 355
rect 296 351 297 355
rect 291 347 297 351
rect 299 352 305 356
rect 299 348 300 352
rect 304 348 305 352
rect 299 347 305 348
rect 424 145 462 146
rect 424 141 432 145
rect 461 141 462 145
rect 424 140 462 141
rect 424 137 462 138
rect 424 133 425 137
rect 454 133 462 137
rect 424 132 462 133
rect 424 129 462 130
rect 424 125 432 129
rect 461 125 462 129
rect 424 124 462 125
rect 424 121 462 122
rect 424 117 425 121
rect 454 117 462 121
rect 424 116 462 117
rect 424 113 462 114
rect 424 109 432 113
rect 461 109 462 113
rect 424 108 462 109
rect 424 105 462 106
rect 424 101 425 105
rect 454 101 462 105
rect 424 100 462 101
rect 424 97 462 98
rect 424 93 432 97
rect 461 93 462 97
rect 424 92 462 93
rect 424 89 462 90
rect 424 85 425 89
rect 454 85 462 89
rect 424 84 462 85
rect 424 81 462 82
rect 424 77 432 81
rect 461 77 462 81
rect 424 76 462 77
rect 424 73 462 74
rect 424 69 425 73
rect 454 69 462 73
rect 424 68 462 69
rect 424 65 462 66
rect 424 61 432 65
rect 461 61 462 65
rect 424 60 462 61
rect 424 57 462 58
rect 424 53 425 57
rect 454 53 462 57
rect 424 52 462 53
rect 424 49 462 50
rect 424 45 432 49
rect 461 45 462 49
rect 424 44 462 45
rect 424 41 462 42
rect 424 37 425 41
rect 454 37 462 41
rect 424 36 462 37
rect 424 33 462 34
rect 424 29 432 33
rect 461 29 462 33
rect 424 28 462 29
rect 424 25 462 26
rect 424 21 425 25
rect 454 21 462 25
rect 424 20 462 21
rect 424 17 462 18
rect 424 13 432 17
rect 461 13 462 17
rect 424 12 462 13
<< pdiffusion >>
rect 124 347 142 348
rect 124 343 125 347
rect 129 343 131 347
rect 135 343 137 347
rect 141 343 142 347
rect 124 341 142 343
rect 124 337 125 341
rect 129 337 131 341
rect 135 337 137 341
rect 141 337 142 341
rect 124 336 142 337
rect 180 347 198 348
rect 180 343 181 347
rect 185 343 187 347
rect 191 343 193 347
rect 197 343 198 347
rect 180 341 198 343
rect 180 337 181 341
rect 185 337 187 341
rect 191 337 193 341
rect 197 337 198 341
rect 180 336 198 337
rect 320 354 326 355
rect 320 350 321 354
rect 325 350 326 354
rect 320 344 326 350
rect 249 334 255 335
rect 249 330 250 334
rect 254 330 255 334
rect 249 328 255 330
rect 249 324 250 328
rect 254 324 255 328
rect 249 322 255 324
rect 249 318 250 322
rect 254 318 255 322
rect 249 317 255 318
rect 257 317 260 335
rect 262 334 268 335
rect 262 330 263 334
rect 267 330 268 334
rect 262 328 268 330
rect 262 324 263 328
rect 267 324 268 328
rect 262 322 268 324
rect 262 318 263 322
rect 267 318 268 322
rect 262 317 268 318
rect 270 317 273 335
rect 275 334 281 335
rect 275 330 276 334
rect 280 330 281 334
rect 275 328 281 330
rect 275 324 276 328
rect 280 324 281 328
rect 275 322 281 324
rect 275 318 276 322
rect 280 318 281 322
rect 275 317 281 318
rect 283 317 289 335
rect 291 334 297 335
rect 291 330 292 334
rect 296 330 297 334
rect 291 328 297 330
rect 291 324 292 328
rect 296 324 297 328
rect 291 322 297 324
rect 291 318 292 322
rect 296 318 297 322
rect 291 317 297 318
rect 299 334 305 335
rect 299 330 300 334
rect 304 330 305 334
rect 299 328 305 330
rect 299 324 300 328
rect 304 324 305 328
rect 299 322 305 324
rect 299 318 300 322
rect 304 318 305 322
rect 299 317 305 318
rect 320 340 321 344
rect 325 340 326 344
rect 320 334 326 340
rect 320 330 321 334
rect 325 330 326 334
rect 320 317 326 330
rect 328 347 334 355
rect 328 318 329 347
rect 333 318 334 347
rect 328 317 334 318
rect 336 354 342 355
rect 336 350 337 354
rect 341 350 342 354
rect 336 344 342 350
rect 336 340 337 344
rect 341 340 342 344
rect 336 334 342 340
rect 336 330 337 334
rect 341 330 342 334
rect 336 317 342 330
rect 344 347 350 355
rect 344 318 345 347
rect 349 318 350 347
rect 344 317 350 318
rect 352 354 358 355
rect 352 350 353 354
rect 357 350 358 354
rect 352 344 358 350
rect 352 340 353 344
rect 357 340 358 344
rect 352 334 358 340
rect 352 330 353 334
rect 357 330 358 334
rect 352 317 358 330
rect 360 347 366 355
rect 360 318 361 347
rect 365 318 366 347
rect 360 317 366 318
rect 368 354 374 355
rect 368 350 369 354
rect 373 350 374 354
rect 368 344 374 350
rect 368 340 369 344
rect 373 340 374 344
rect 368 334 374 340
rect 368 330 369 334
rect 373 330 374 334
rect 368 317 374 330
rect 376 347 382 355
rect 376 318 377 347
rect 381 318 382 347
rect 376 317 382 318
rect 384 354 390 355
rect 384 350 385 354
rect 389 350 390 354
rect 384 344 390 350
rect 384 340 385 344
rect 389 340 390 344
rect 384 334 390 340
rect 384 330 385 334
rect 389 330 390 334
rect 384 317 390 330
rect 392 347 398 355
rect 392 318 393 347
rect 397 318 398 347
rect 392 317 398 318
rect 400 354 406 355
rect 400 350 401 354
rect 405 350 406 354
rect 400 344 406 350
rect 400 340 401 344
rect 405 340 406 344
rect 400 334 406 340
rect 400 330 401 334
rect 405 330 406 334
rect 400 317 406 330
rect 408 347 414 355
rect 408 318 409 347
rect 413 318 414 347
rect 408 317 414 318
rect 416 354 422 355
rect 416 350 417 354
rect 421 350 422 354
rect 416 344 422 350
rect 416 340 417 344
rect 421 340 422 344
rect 416 334 422 340
rect 416 330 417 334
rect 421 330 422 334
rect 416 317 422 330
rect 424 347 430 355
rect 424 318 425 347
rect 429 318 430 347
rect 424 317 430 318
rect 432 354 438 355
rect 432 350 433 354
rect 437 350 438 354
rect 432 344 438 350
rect 432 340 433 344
rect 437 340 438 344
rect 432 334 438 340
rect 432 330 433 334
rect 437 330 438 334
rect 432 317 438 330
rect 440 347 446 355
rect 440 318 441 347
rect 445 318 446 347
rect 440 317 446 318
rect 448 354 454 355
rect 448 350 449 354
rect 453 350 454 354
rect 448 344 454 350
rect 448 340 449 344
rect 453 340 454 344
rect 448 334 454 340
rect 448 330 449 334
rect 453 330 454 334
rect 448 317 454 330
rect 424 301 462 302
rect 424 297 434 301
rect 438 297 444 301
rect 448 297 454 301
rect 458 297 462 301
rect 424 296 462 297
rect 424 293 462 294
rect 424 289 425 293
rect 454 289 462 293
rect 424 288 462 289
rect 424 285 462 286
rect 424 281 434 285
rect 438 281 444 285
rect 448 281 454 285
rect 458 281 462 285
rect 424 280 462 281
rect 424 277 462 278
rect 424 273 425 277
rect 454 273 462 277
rect 424 272 462 273
rect 424 269 462 270
rect 424 265 434 269
rect 438 265 444 269
rect 448 265 454 269
rect 458 265 462 269
rect 424 264 462 265
rect 424 261 462 262
rect 424 257 425 261
rect 454 257 462 261
rect 424 256 462 257
rect 424 253 462 254
rect 424 249 434 253
rect 438 249 444 253
rect 448 249 454 253
rect 458 249 462 253
rect 424 248 462 249
rect 424 245 462 246
rect 424 241 425 245
rect 454 241 462 245
rect 424 240 462 241
rect 424 237 462 238
rect 424 233 434 237
rect 438 233 444 237
rect 448 233 454 237
rect 458 233 462 237
rect 424 232 462 233
rect 424 229 462 230
rect 424 225 425 229
rect 454 225 462 229
rect 424 224 462 225
rect 424 221 462 222
rect 424 217 434 221
rect 438 217 444 221
rect 448 217 454 221
rect 458 217 462 221
rect 424 216 462 217
rect 424 213 462 214
rect 424 209 425 213
rect 454 209 462 213
rect 424 208 462 209
rect 424 205 462 206
rect 424 201 434 205
rect 438 201 444 205
rect 448 201 454 205
rect 458 201 462 205
rect 424 200 462 201
rect 424 197 462 198
rect 424 193 425 197
rect 454 193 462 197
rect 424 192 462 193
rect 424 189 462 190
rect 424 185 434 189
rect 438 185 444 189
rect 448 185 454 189
rect 458 185 462 189
rect 424 184 462 185
rect 424 181 462 182
rect 424 177 425 181
rect 454 177 462 181
rect 424 176 462 177
rect 424 173 462 174
rect 424 169 434 173
rect 438 169 444 173
rect 448 169 454 173
rect 458 169 462 173
rect 424 168 462 169
<< ndcontact >>
rect 35 355 39 359
rect 41 355 45 359
rect 35 349 39 353
rect 41 349 45 353
rect 35 343 39 347
rect 41 343 45 347
rect 35 337 39 341
rect 41 337 45 341
rect 35 331 39 335
rect 41 331 45 335
rect 35 325 39 329
rect 41 325 45 329
rect 61 355 65 359
rect 67 355 71 359
rect 61 349 65 353
rect 67 349 71 353
rect 61 343 65 347
rect 67 343 71 347
rect 61 337 65 341
rect 67 337 71 341
rect 61 331 65 335
rect 67 331 71 335
rect 61 325 65 329
rect 67 325 71 329
rect 87 355 91 359
rect 93 355 97 359
rect 87 349 91 353
rect 93 349 97 353
rect 87 343 91 347
rect 93 343 97 347
rect 87 337 91 341
rect 93 337 97 341
rect 87 331 91 335
rect 93 331 97 335
rect 87 325 91 329
rect 93 325 97 329
rect 250 351 254 355
rect 263 348 267 352
rect 276 351 280 355
rect 284 348 288 352
rect 292 351 296 355
rect 300 348 304 352
rect 432 141 461 145
rect 425 133 454 137
rect 432 125 461 129
rect 425 117 454 121
rect 432 109 461 113
rect 425 101 454 105
rect 432 93 461 97
rect 425 85 454 89
rect 432 77 461 81
rect 425 69 454 73
rect 432 61 461 65
rect 425 53 454 57
rect 432 45 461 49
rect 425 37 454 41
rect 432 29 461 33
rect 425 21 454 25
rect 432 13 461 17
<< pdcontact >>
rect 125 343 129 347
rect 131 343 135 347
rect 137 343 141 347
rect 125 337 129 341
rect 131 337 135 341
rect 137 337 141 341
rect 181 343 185 347
rect 187 343 191 347
rect 193 343 197 347
rect 181 337 185 341
rect 187 337 191 341
rect 193 337 197 341
rect 321 350 325 354
rect 250 330 254 334
rect 250 324 254 328
rect 250 318 254 322
rect 263 330 267 334
rect 263 324 267 328
rect 263 318 267 322
rect 276 330 280 334
rect 276 324 280 328
rect 276 318 280 322
rect 292 330 296 334
rect 292 324 296 328
rect 292 318 296 322
rect 300 330 304 334
rect 300 324 304 328
rect 300 318 304 322
rect 321 340 325 344
rect 321 330 325 334
rect 329 318 333 347
rect 337 350 341 354
rect 337 340 341 344
rect 337 330 341 334
rect 345 318 349 347
rect 353 350 357 354
rect 353 340 357 344
rect 353 330 357 334
rect 361 318 365 347
rect 369 350 373 354
rect 369 340 373 344
rect 369 330 373 334
rect 377 318 381 347
rect 385 350 389 354
rect 385 340 389 344
rect 385 330 389 334
rect 393 318 397 347
rect 401 350 405 354
rect 401 340 405 344
rect 401 330 405 334
rect 409 318 413 347
rect 417 350 421 354
rect 417 340 421 344
rect 417 330 421 334
rect 425 318 429 347
rect 433 350 437 354
rect 433 340 437 344
rect 433 330 437 334
rect 441 318 445 347
rect 449 350 453 354
rect 449 340 453 344
rect 449 330 453 334
rect 434 297 438 301
rect 444 297 448 301
rect 454 297 458 301
rect 425 289 454 293
rect 434 281 438 285
rect 444 281 448 285
rect 454 281 458 285
rect 425 273 454 277
rect 434 265 438 269
rect 444 265 448 269
rect 454 265 458 269
rect 425 257 454 261
rect 434 249 438 253
rect 444 249 448 253
rect 454 249 458 253
rect 425 241 454 245
rect 434 233 438 237
rect 444 233 448 237
rect 454 233 458 237
rect 425 225 454 229
rect 434 217 438 221
rect 444 217 448 221
rect 454 217 458 221
rect 425 209 454 213
rect 434 201 438 205
rect 444 201 448 205
rect 454 201 458 205
rect 425 193 454 197
rect 434 185 438 189
rect 444 185 448 189
rect 454 185 458 189
rect 425 177 454 181
rect 434 169 438 173
rect 444 169 448 173
rect 454 169 458 173
<< psubstratepdiff >>
rect 24 361 30 364
rect 24 357 25 361
rect 29 357 30 361
rect 50 361 56 364
rect 24 355 30 357
rect 24 351 25 355
rect 29 351 30 355
rect 24 349 30 351
rect 24 345 25 349
rect 29 345 30 349
rect 24 343 30 345
rect 24 339 25 343
rect 29 339 30 343
rect 24 337 30 339
rect 24 333 25 337
rect 29 333 30 337
rect 24 331 30 333
rect 24 327 25 331
rect 29 327 30 331
rect 24 320 30 327
rect 50 357 51 361
rect 55 357 56 361
rect 76 361 82 364
rect 50 355 56 357
rect 50 351 51 355
rect 55 351 56 355
rect 50 349 56 351
rect 50 345 51 349
rect 55 345 56 349
rect 50 343 56 345
rect 50 339 51 343
rect 55 339 56 343
rect 50 337 56 339
rect 50 333 51 337
rect 55 333 56 337
rect 50 331 56 333
rect 50 327 51 331
rect 55 327 56 331
rect 50 320 56 327
rect 76 357 77 361
rect 81 357 82 361
rect 102 361 108 364
rect 76 355 82 357
rect 76 351 77 355
rect 81 351 82 355
rect 76 349 82 351
rect 76 345 77 349
rect 81 345 82 349
rect 76 343 82 345
rect 76 339 77 343
rect 81 339 82 343
rect 76 337 82 339
rect 76 333 77 337
rect 81 333 82 337
rect 76 331 82 333
rect 76 327 77 331
rect 81 327 82 331
rect 76 320 82 327
rect 102 357 103 361
rect 107 357 108 361
rect 158 361 164 364
rect 102 355 108 357
rect 102 351 103 355
rect 107 351 108 355
rect 102 349 108 351
rect 102 345 103 349
rect 107 345 108 349
rect 102 343 108 345
rect 102 339 103 343
rect 107 339 108 343
rect 102 337 108 339
rect 102 333 103 337
rect 107 333 108 337
rect 102 331 108 333
rect 102 327 103 331
rect 107 327 108 331
rect 102 320 108 327
rect 158 357 159 361
rect 163 357 164 361
rect 214 361 220 364
rect 158 355 164 357
rect 158 351 159 355
rect 163 351 164 355
rect 158 349 164 351
rect 158 345 159 349
rect 163 345 164 349
rect 158 343 164 345
rect 158 339 159 343
rect 163 339 164 343
rect 158 337 164 339
rect 158 333 159 337
rect 163 333 164 337
rect 158 331 164 333
rect 158 327 159 331
rect 163 327 164 331
rect 158 320 164 327
rect 214 357 215 361
rect 219 357 220 361
rect 214 355 220 357
rect 214 351 215 355
rect 219 351 220 355
rect 214 349 220 351
rect 214 345 215 349
rect 219 345 220 349
rect 214 343 220 345
rect 214 339 215 343
rect 219 339 220 343
rect 214 337 220 339
rect 214 333 215 337
rect 219 333 220 337
rect 214 331 220 333
rect 214 327 215 331
rect 219 327 220 331
rect 214 320 220 327
rect 24 314 220 320
rect 424 151 462 152
rect 424 147 432 151
rect 461 147 462 151
rect 424 146 462 147
rect 424 11 462 12
rect 424 7 432 11
rect 461 7 462 11
rect 424 6 462 7
<< nsubstratendiff >>
rect 114 357 152 358
rect 114 353 115 357
rect 119 353 127 357
rect 131 353 135 357
rect 139 353 147 357
rect 151 353 152 357
rect 114 352 152 353
rect 114 349 120 352
rect 114 345 115 349
rect 119 345 120 349
rect 146 349 152 352
rect 114 341 120 345
rect 114 337 115 341
rect 119 337 120 341
rect 114 333 120 337
rect 146 345 147 349
rect 151 345 152 349
rect 146 341 152 345
rect 146 337 147 341
rect 151 337 152 341
rect 114 329 115 333
rect 119 332 120 333
rect 146 333 152 337
rect 146 332 147 333
rect 119 329 147 332
rect 151 329 152 333
rect 114 326 152 329
rect 170 357 208 358
rect 170 353 171 357
rect 175 353 183 357
rect 187 353 191 357
rect 195 353 203 357
rect 207 353 208 357
rect 170 352 208 353
rect 170 349 176 352
rect 170 345 171 349
rect 175 345 176 349
rect 202 349 208 352
rect 170 341 176 345
rect 170 337 171 341
rect 175 337 176 341
rect 170 333 176 337
rect 202 345 203 349
rect 207 345 208 349
rect 202 341 208 345
rect 202 337 203 341
rect 207 337 208 341
rect 170 329 171 333
rect 175 332 176 333
rect 202 333 208 337
rect 202 332 203 333
rect 175 329 203 332
rect 207 329 208 333
rect 170 326 208 329
rect 314 354 320 355
rect 314 350 315 354
rect 319 350 320 354
rect 314 344 320 350
rect 314 340 315 344
rect 319 340 320 344
rect 314 334 320 340
rect 314 330 315 334
rect 319 330 320 334
rect 314 317 320 330
rect 454 349 460 355
rect 454 345 455 349
rect 459 345 460 349
rect 454 339 460 345
rect 454 335 455 339
rect 459 335 460 339
rect 454 329 460 335
rect 454 325 455 329
rect 459 325 460 329
rect 454 317 460 325
rect 424 307 462 308
rect 424 303 429 307
rect 433 303 439 307
rect 443 303 449 307
rect 453 303 462 307
rect 424 302 462 303
rect 424 167 462 168
rect 424 163 429 167
rect 433 163 439 167
rect 443 163 449 167
rect 453 163 462 167
rect 424 162 462 163
<< psubstratepcontact >>
rect 25 357 29 361
rect 25 351 29 355
rect 25 345 29 349
rect 25 339 29 343
rect 25 333 29 337
rect 25 327 29 331
rect 51 357 55 361
rect 51 351 55 355
rect 51 345 55 349
rect 51 339 55 343
rect 51 333 55 337
rect 51 327 55 331
rect 77 357 81 361
rect 77 351 81 355
rect 77 345 81 349
rect 77 339 81 343
rect 77 333 81 337
rect 77 327 81 331
rect 103 357 107 361
rect 103 351 107 355
rect 103 345 107 349
rect 103 339 107 343
rect 103 333 107 337
rect 103 327 107 331
rect 159 357 163 361
rect 159 351 163 355
rect 159 345 163 349
rect 159 339 163 343
rect 159 333 163 337
rect 159 327 163 331
rect 215 357 219 361
rect 215 351 219 355
rect 215 345 219 349
rect 215 339 219 343
rect 215 333 219 337
rect 215 327 219 331
rect 432 147 461 151
rect 432 7 461 11
<< nsubstratencontact >>
rect 115 353 119 357
rect 127 353 131 357
rect 135 353 139 357
rect 147 353 151 357
rect 115 345 119 349
rect 115 337 119 341
rect 147 345 151 349
rect 147 337 151 341
rect 115 329 119 333
rect 147 329 151 333
rect 171 353 175 357
rect 183 353 187 357
rect 191 353 195 357
rect 203 353 207 357
rect 171 345 175 349
rect 171 337 175 341
rect 203 345 207 349
rect 203 337 207 341
rect 171 329 175 333
rect 203 329 207 333
rect 315 350 319 354
rect 315 340 319 344
rect 315 330 319 334
rect 455 345 459 349
rect 455 335 459 339
rect 455 325 459 329
rect 429 303 433 307
rect 439 303 443 307
rect 449 303 453 307
rect 429 163 433 167
rect 439 163 443 167
rect 449 163 453 167
<< polysilicon >>
rect 9 357 21 358
rect 9 343 10 357
rect 14 343 16 357
rect 20 343 21 357
rect 9 25 21 343
rect 241 362 299 363
rect 241 358 242 362
rect 246 361 299 362
rect 246 358 247 361
rect 241 357 247 358
rect 255 356 257 361
rect 260 356 262 358
rect 268 356 270 358
rect 273 356 275 361
rect 281 356 283 358
rect 289 356 291 358
rect 297 356 299 361
rect 311 362 470 363
rect 311 358 317 362
rect 321 358 327 362
rect 331 358 470 362
rect 311 357 470 358
rect 326 355 328 357
rect 334 355 336 357
rect 342 355 344 357
rect 350 355 352 357
rect 358 355 360 357
rect 366 355 368 357
rect 374 355 376 357
rect 382 355 384 357
rect 390 355 392 357
rect 398 355 400 357
rect 406 355 408 357
rect 414 355 416 357
rect 422 355 424 357
rect 430 355 432 357
rect 438 355 440 357
rect 446 355 448 357
rect 255 335 257 347
rect 260 342 262 347
rect 268 342 270 347
rect 273 345 275 347
rect 281 342 283 347
rect 260 340 283 342
rect 260 335 262 340
rect 268 335 270 337
rect 273 335 275 340
rect 281 335 283 340
rect 289 335 291 347
rect 297 335 299 347
rect 302 343 308 344
rect 302 339 303 343
rect 307 339 308 343
rect 302 338 308 339
rect 234 315 240 316
rect 255 315 257 317
rect 24 301 51 313
rect 234 311 235 315
rect 239 312 240 315
rect 260 312 262 317
rect 239 311 262 312
rect 234 310 262 311
rect 268 312 270 317
rect 273 315 275 317
rect 281 315 283 317
rect 289 312 291 317
rect 297 315 299 317
rect 306 312 308 338
rect 326 315 328 317
rect 334 315 336 317
rect 342 315 344 317
rect 350 315 352 317
rect 358 315 360 317
rect 366 315 368 317
rect 374 315 376 317
rect 382 315 384 317
rect 390 315 392 317
rect 398 315 400 317
rect 406 315 408 317
rect 414 315 416 317
rect 422 315 424 317
rect 430 315 432 317
rect 438 315 440 317
rect 446 315 448 317
rect 268 310 308 312
rect 24 25 36 301
rect 9 13 36 25
rect 39 31 51 301
rect 464 296 470 357
rect 422 294 424 296
rect 462 294 470 296
rect 464 288 470 294
rect 422 286 424 288
rect 462 286 470 288
rect 464 280 470 286
rect 422 278 424 280
rect 462 278 470 280
rect 464 272 470 278
rect 422 270 424 272
rect 462 270 470 272
rect 464 264 470 270
rect 422 262 424 264
rect 462 262 470 264
rect 464 256 470 262
rect 422 254 424 256
rect 462 254 470 256
rect 464 248 470 254
rect 422 246 424 248
rect 462 246 470 248
rect 464 240 470 246
rect 422 238 424 240
rect 462 238 470 240
rect 464 232 470 238
rect 422 230 424 232
rect 462 230 470 232
rect 464 224 470 230
rect 422 222 424 224
rect 462 222 470 224
rect 464 216 470 222
rect 422 214 424 216
rect 462 214 470 216
rect 464 208 470 214
rect 422 206 424 208
rect 462 206 470 208
rect 464 200 470 206
rect 422 198 424 200
rect 462 198 470 200
rect 464 192 470 198
rect 422 190 424 192
rect 462 190 470 192
rect 464 184 470 190
rect 422 182 424 184
rect 462 182 470 184
rect 464 176 470 182
rect 422 174 424 176
rect 462 174 470 176
rect 433 158 470 159
rect 433 154 439 158
rect 443 154 449 158
rect 453 154 470 158
rect 433 153 470 154
rect 464 140 470 153
rect 422 138 424 140
rect 462 138 470 140
rect 464 132 470 138
rect 422 130 424 132
rect 462 130 470 132
rect 464 124 470 130
rect 422 122 424 124
rect 462 122 470 124
rect 464 116 470 122
rect 422 114 424 116
rect 462 114 470 116
rect 464 108 470 114
rect 422 106 424 108
rect 462 106 470 108
rect 464 100 470 106
rect 422 98 424 100
rect 462 98 470 100
rect 464 92 470 98
rect 422 90 424 92
rect 462 90 470 92
rect 464 84 470 90
rect 422 82 424 84
rect 462 82 470 84
rect 464 76 470 82
rect 422 74 424 76
rect 462 74 470 76
rect 464 68 470 74
rect 422 66 424 68
rect 462 66 470 68
rect 464 60 470 66
rect 422 58 424 60
rect 462 58 470 60
rect 464 52 470 58
rect 422 50 424 52
rect 462 50 470 52
rect 464 44 470 50
rect 422 42 424 44
rect 462 42 470 44
rect 464 36 470 42
rect 422 34 424 36
rect 462 34 470 36
rect 39 29 52 31
rect 39 15 41 29
rect 50 15 52 29
rect 464 28 470 34
rect 422 26 424 28
rect 462 26 470 28
rect 464 20 470 26
rect 422 18 424 20
rect 462 18 470 20
rect 39 13 52 15
<< polycontact >>
rect 10 343 14 357
rect 16 343 20 357
rect 242 358 246 362
rect 317 358 321 362
rect 327 358 331 362
rect 303 339 307 343
rect 235 311 239 315
rect 439 154 443 158
rect 449 154 453 158
rect 41 15 50 29
<< metal1 >>
rect -2 365 224 369
rect -2 3 2 365
rect 25 361 29 365
rect 9 357 21 358
rect 9 343 10 357
rect 14 343 16 357
rect 20 343 21 357
rect 9 323 21 343
rect 51 361 55 365
rect 25 355 29 357
rect 25 349 29 351
rect 25 343 29 345
rect 25 337 29 339
rect 25 331 29 333
rect 39 355 41 359
rect 35 353 45 355
rect 39 349 41 353
rect 35 347 45 349
rect 39 343 41 347
rect 35 341 45 343
rect 39 337 41 341
rect 35 335 45 337
rect 39 331 41 335
rect 35 329 45 331
rect 39 325 41 329
rect 77 361 81 365
rect 51 355 55 357
rect 51 349 55 351
rect 51 343 55 345
rect 51 337 55 339
rect 51 331 55 333
rect 65 355 67 359
rect 61 353 71 355
rect 65 349 67 353
rect 61 347 71 349
rect 65 343 67 347
rect 61 341 71 343
rect 65 337 67 341
rect 61 335 71 337
rect 65 331 67 335
rect 61 329 71 331
rect 35 323 45 325
rect 65 325 67 329
rect 103 361 107 365
rect 77 355 81 357
rect 77 349 81 351
rect 77 343 81 345
rect 77 337 81 339
rect 77 331 81 333
rect 91 355 93 359
rect 87 353 97 355
rect 91 349 93 353
rect 87 347 97 349
rect 91 343 93 347
rect 87 341 97 343
rect 91 337 93 341
rect 87 335 97 337
rect 91 331 93 335
rect 87 329 97 331
rect 61 323 71 325
rect 91 325 93 329
rect 159 361 163 365
rect 215 361 219 365
rect 103 355 107 357
rect 103 349 107 351
rect 103 343 107 345
rect 103 337 107 339
rect 103 331 107 333
rect 119 353 123 357
rect 143 353 147 357
rect 129 343 131 347
rect 135 343 137 347
rect 125 341 141 343
rect 129 337 131 341
rect 135 337 137 341
rect 87 323 97 325
rect 125 323 141 337
rect 159 355 163 357
rect 159 349 163 351
rect 159 343 163 345
rect 159 337 163 339
rect 159 331 163 333
rect 175 353 179 357
rect 199 353 203 357
rect 185 343 187 347
rect 191 343 193 347
rect 181 341 197 343
rect 185 337 187 341
rect 191 337 193 341
rect 181 323 197 337
rect 215 355 219 357
rect 215 349 219 351
rect 215 343 219 345
rect 215 337 219 339
rect 215 331 219 333
rect 229 323 232 513
rect 9 310 232 323
rect 235 315 239 513
rect 242 362 245 513
rect 250 365 476 369
rect 250 355 254 365
rect 276 355 280 365
rect 292 355 296 365
rect 316 358 317 362
rect 321 358 322 362
rect 326 358 327 362
rect 263 346 267 348
rect 254 342 267 346
rect 284 346 288 348
rect 250 340 254 342
rect 284 340 288 342
rect 250 334 254 336
rect 276 336 284 340
rect 300 343 304 348
rect 319 350 321 354
rect 315 349 325 350
rect 319 345 321 349
rect 337 349 341 350
rect 315 344 325 345
rect 300 339 303 343
rect 319 340 321 344
rect 315 339 325 340
rect 276 334 280 336
rect 300 334 304 339
rect 250 328 254 330
rect 250 322 254 324
rect 263 328 267 330
rect 263 322 267 324
rect 276 328 280 330
rect 276 322 280 324
rect 292 328 296 330
rect 292 322 296 324
rect 300 328 304 330
rect 300 322 304 324
rect 319 335 321 339
rect 315 334 325 335
rect 319 330 321 334
rect 315 329 325 330
rect 319 325 321 329
rect 263 314 267 318
rect 292 314 296 318
rect 315 314 325 325
rect 263 310 325 314
rect 353 349 357 350
rect 337 344 341 345
rect 337 339 341 340
rect 337 334 341 335
rect 337 329 341 330
rect 333 318 345 322
rect 369 349 373 350
rect 353 344 357 345
rect 353 339 357 340
rect 353 334 357 335
rect 353 329 357 330
rect 349 318 361 322
rect 385 349 389 350
rect 369 344 373 345
rect 369 339 373 340
rect 369 334 373 335
rect 369 329 373 330
rect 365 318 377 322
rect 401 349 405 350
rect 385 344 389 345
rect 385 339 389 340
rect 385 334 389 335
rect 385 329 389 330
rect 381 318 393 322
rect 417 349 421 350
rect 401 344 405 345
rect 401 339 405 340
rect 401 334 405 335
rect 401 329 405 330
rect 397 318 409 322
rect 433 349 437 350
rect 417 344 421 345
rect 417 339 421 340
rect 417 334 421 335
rect 417 329 421 330
rect 413 318 425 322
rect 453 350 455 354
rect 449 349 459 350
rect 433 344 437 345
rect 433 339 437 340
rect 433 334 437 335
rect 433 329 437 330
rect 429 318 441 322
rect 453 345 455 349
rect 449 344 459 345
rect 453 340 455 344
rect 449 339 459 340
rect 453 335 455 339
rect 449 334 459 335
rect 453 330 455 334
rect 449 329 459 330
rect 453 325 455 329
rect 329 310 445 318
rect 39 29 107 31
rect 39 15 41 29
rect 50 15 107 29
rect 39 13 107 15
rect 329 0 425 310
rect 433 303 434 307
rect 438 303 439 307
rect 443 303 444 307
rect 448 303 449 307
rect 453 303 454 307
rect 429 301 458 303
rect 433 297 434 301
rect 438 297 439 301
rect 443 297 444 301
rect 448 297 449 301
rect 453 297 454 301
rect 433 281 434 285
rect 438 281 439 285
rect 443 281 444 285
rect 448 281 449 285
rect 453 281 454 285
rect 433 265 434 269
rect 438 265 439 269
rect 443 265 444 269
rect 448 265 449 269
rect 453 265 454 269
rect 433 249 434 253
rect 438 249 439 253
rect 443 249 444 253
rect 448 249 449 253
rect 453 249 454 253
rect 433 233 434 237
rect 438 233 439 237
rect 443 233 444 237
rect 448 233 449 237
rect 453 233 454 237
rect 433 217 434 221
rect 438 217 439 221
rect 443 217 444 221
rect 448 217 449 221
rect 453 217 454 221
rect 433 201 434 205
rect 438 201 439 205
rect 443 201 444 205
rect 448 201 449 205
rect 453 201 454 205
rect 433 185 434 189
rect 438 185 439 189
rect 443 185 444 189
rect 448 185 449 189
rect 453 185 454 189
rect 433 169 434 173
rect 438 169 439 173
rect 443 169 444 173
rect 448 169 449 173
rect 453 169 454 173
rect 429 167 458 169
rect 433 163 434 167
rect 438 163 439 167
rect 443 163 444 167
rect 448 163 449 167
rect 453 163 454 167
rect 438 154 439 158
rect 443 154 444 158
rect 448 154 449 158
rect 462 151 476 365
rect 461 147 476 151
rect 432 145 476 147
rect 461 141 476 145
rect 462 129 476 141
rect 461 125 476 129
rect 462 113 476 125
rect 461 109 476 113
rect 462 97 476 109
rect 461 93 476 97
rect 462 81 476 93
rect 461 77 476 81
rect 462 65 476 77
rect 461 61 476 65
rect 462 49 476 61
rect 461 45 476 49
rect 462 33 476 45
rect 461 29 476 33
rect 462 17 476 29
rect 461 13 476 17
rect 432 11 476 13
rect 461 7 476 11
rect 462 3 476 7
<< m2contact >>
rect 123 353 127 357
rect 131 353 135 357
rect 139 353 143 357
rect 115 349 119 353
rect 147 349 151 353
rect 115 341 119 345
rect 115 333 119 337
rect 147 341 151 345
rect 147 333 151 337
rect 179 353 183 357
rect 187 353 191 357
rect 195 353 199 357
rect 171 349 175 353
rect 203 349 207 353
rect 171 341 175 345
rect 171 333 175 337
rect 203 341 207 345
rect 203 333 207 337
rect 312 358 316 362
rect 322 358 326 362
rect 250 342 254 346
rect 284 342 288 346
rect 250 336 254 340
rect 284 336 288 340
rect 315 345 319 349
rect 321 345 325 349
rect 315 335 319 339
rect 321 335 325 339
rect 315 325 319 329
rect 321 325 325 329
rect 337 345 341 349
rect 337 335 341 339
rect 337 325 341 329
rect 353 345 357 349
rect 353 335 357 339
rect 353 325 357 329
rect 369 345 373 349
rect 369 335 373 339
rect 369 325 373 329
rect 385 345 389 349
rect 385 335 389 339
rect 385 325 389 329
rect 401 345 405 349
rect 401 335 405 339
rect 401 325 405 329
rect 417 345 421 349
rect 417 335 421 339
rect 417 325 421 329
rect 433 345 437 349
rect 455 350 459 354
rect 433 335 437 339
rect 433 325 437 329
rect 449 345 453 349
rect 455 340 459 344
rect 449 335 453 339
rect 455 330 459 334
rect 449 325 453 329
rect 434 303 438 307
rect 444 303 448 307
rect 454 303 458 307
rect 429 297 433 301
rect 439 297 443 301
rect 449 297 453 301
rect 429 281 433 285
rect 439 281 443 285
rect 449 281 453 285
rect 429 265 433 269
rect 439 265 443 269
rect 449 265 453 269
rect 429 249 433 253
rect 439 249 443 253
rect 449 249 453 253
rect 429 233 433 237
rect 439 233 443 237
rect 449 233 453 237
rect 429 217 433 221
rect 439 217 443 221
rect 449 217 453 221
rect 429 201 433 205
rect 439 201 443 205
rect 449 201 453 205
rect 429 185 433 189
rect 439 185 443 189
rect 449 185 453 189
rect 429 169 433 173
rect 439 169 443 173
rect 449 169 453 173
rect 434 163 438 167
rect 444 163 448 167
rect 454 163 458 167
rect 434 154 438 158
rect 444 154 448 158
<< metal2 >>
rect 114 357 152 367
rect 114 353 123 357
rect 127 353 131 357
rect 135 353 139 357
rect 143 353 152 357
rect 114 349 115 353
rect 119 352 147 353
rect 119 349 120 352
rect 114 345 120 349
rect 114 341 115 345
rect 119 341 120 345
rect 114 337 120 341
rect 114 333 115 337
rect 119 333 120 337
rect 114 332 120 333
rect 146 349 147 352
rect 151 349 152 353
rect 146 345 152 349
rect 146 341 147 345
rect 151 341 152 345
rect 146 337 152 341
rect 146 333 147 337
rect 151 333 152 337
rect 146 332 152 333
rect 170 357 208 367
rect 170 353 179 357
rect 183 353 187 357
rect 191 353 195 357
rect 199 353 208 357
rect 170 349 171 353
rect 175 352 203 353
rect 175 349 176 352
rect 170 345 176 349
rect 170 341 171 345
rect 175 341 176 345
rect 170 337 176 341
rect 170 333 171 337
rect 175 333 176 337
rect 170 332 176 333
rect 202 349 203 352
rect 207 349 208 353
rect 202 345 208 349
rect 202 341 203 345
rect 207 341 208 345
rect 202 337 208 341
rect 202 333 203 337
rect 207 333 208 337
rect 250 358 312 362
rect 316 358 322 362
rect 250 346 254 358
rect 337 354 459 367
rect 337 350 455 354
rect 337 349 459 350
rect 250 340 254 342
rect 284 340 288 342
rect 202 332 208 333
rect 284 314 288 336
rect 319 345 321 349
rect 325 345 337 349
rect 341 345 353 349
rect 357 345 369 349
rect 373 345 385 349
rect 389 345 401 349
rect 405 345 417 349
rect 421 345 433 349
rect 437 345 449 349
rect 453 345 459 349
rect 315 344 459 345
rect 315 340 455 344
rect 315 339 459 340
rect 319 335 321 339
rect 325 335 337 339
rect 341 335 353 339
rect 357 335 369 339
rect 373 335 385 339
rect 389 335 401 339
rect 405 335 417 339
rect 421 335 433 339
rect 437 335 449 339
rect 453 335 459 339
rect 315 334 459 335
rect 315 330 455 334
rect 315 329 459 330
rect 319 325 321 329
rect 325 325 337 329
rect 341 325 353 329
rect 357 325 369 329
rect 373 325 385 329
rect 389 325 401 329
rect 405 325 417 329
rect 421 325 433 329
rect 437 325 449 329
rect 453 325 459 329
rect 284 310 421 314
rect 417 158 421 310
rect 429 307 459 325
rect 429 303 434 307
rect 438 303 444 307
rect 448 303 454 307
rect 458 303 459 307
rect 429 301 459 303
rect 433 297 439 301
rect 443 297 449 301
rect 453 297 459 301
rect 429 285 459 297
rect 433 281 439 285
rect 443 281 449 285
rect 453 281 459 285
rect 429 269 459 281
rect 433 265 439 269
rect 443 265 449 269
rect 453 265 459 269
rect 429 253 459 265
rect 433 249 439 253
rect 443 249 449 253
rect 453 249 459 253
rect 429 237 459 249
rect 433 233 439 237
rect 443 233 449 237
rect 453 233 459 237
rect 429 221 459 233
rect 433 217 439 221
rect 443 217 449 221
rect 453 217 459 221
rect 429 205 459 217
rect 433 201 439 205
rect 443 201 449 205
rect 453 201 459 205
rect 429 189 459 201
rect 433 185 439 189
rect 443 185 449 189
rect 453 185 459 189
rect 429 173 459 185
rect 433 169 439 173
rect 443 169 449 173
rect 453 169 459 173
rect 429 167 459 169
rect 429 163 434 167
rect 438 163 444 167
rect 448 163 454 167
rect 458 163 459 167
rect 417 154 434 158
rect 438 154 444 158
use bondingpad  bondingpad_0
timestamp 1259953556
transform 1 0 107 0 1 0
box 0 0 260 260
<< labels >>
rlabel metal1 237 512 237 512 6 Out
rlabel metal1 244 512 244 512 6 Out_Ena
rlabel metal1 230 512 230 512 6 In
<< end >>
