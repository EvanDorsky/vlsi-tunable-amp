magic
tech scmos
magscale 1 3
timestamp 1419146600
<< metal3 >>
rect 2674 7231 2724 7241
rect 2644 7221 2754 7231
rect 2634 7211 2764 7221
rect 2604 7191 2764 7211
rect 2924 7191 2994 7211
rect 2584 7181 2764 7191
rect 2914 7181 2994 7191
rect 2564 7171 2754 7181
rect 2914 7171 3004 7181
rect 3024 7171 3044 7181
rect 3064 7171 3144 7181
rect 2554 7161 2734 7171
rect 2904 7161 3194 7171
rect 2534 7151 2734 7161
rect 2894 7151 3224 7161
rect 2524 7141 2714 7151
rect 2894 7141 3244 7151
rect 2494 7131 2724 7141
rect 2794 7131 2824 7141
rect 2834 7131 2854 7141
rect 2894 7131 3284 7141
rect 2484 7121 2734 7131
rect 2794 7121 2874 7131
rect 2934 7121 3294 7131
rect 2464 7111 2744 7121
rect 2774 7111 2904 7121
rect 2944 7111 3324 7121
rect 2424 7101 2914 7111
rect 2944 7101 3344 7111
rect 2414 7091 2924 7101
rect 2934 7091 2994 7101
rect 3064 7091 3084 7101
rect 3214 7091 3324 7101
rect 2394 7081 2984 7091
rect 3244 7081 3264 7091
rect 2364 7071 2974 7081
rect 2334 7061 2984 7071
rect 2314 7051 3004 7061
rect 2294 7041 3014 7051
rect 2284 7031 3014 7041
rect 2274 7021 2954 7031
rect 2974 7021 3004 7031
rect 2254 7011 2954 7021
rect 2244 7001 2954 7011
rect 2234 6991 2974 7001
rect 2224 6981 2964 6991
rect 2214 6961 2964 6981
rect 2204 6951 2964 6961
rect 2204 6941 2954 6951
rect 2194 6931 2944 6941
rect 3164 6931 3174 6951
rect 2184 6921 2784 6931
rect 2874 6921 2954 6931
rect 2164 6911 2794 6921
rect 2894 6911 2904 6921
rect 2924 6911 2944 6921
rect 2154 6901 2804 6911
rect 2154 6891 2734 6901
rect 2754 6891 2764 6901
rect 2774 6891 2804 6901
rect 3164 6901 3224 6911
rect 3164 6891 3254 6901
rect 2134 6881 2694 6891
rect 3174 6881 3314 6891
rect 2134 6871 2684 6881
rect 3204 6871 3324 6881
rect 2114 6861 2694 6871
rect 3244 6861 3354 6871
rect 2094 6851 2714 6861
rect 3284 6851 3364 6861
rect 2074 6841 2734 6851
rect 3304 6841 3374 6851
rect 2054 6831 2734 6841
rect 3334 6831 3354 6841
rect 2044 6821 2764 6831
rect 2024 6811 2784 6821
rect 2014 6801 2544 6811
rect 2634 6801 2794 6811
rect 1994 6791 2544 6801
rect 2644 6791 2804 6801
rect 1994 6781 2584 6791
rect 2654 6781 2844 6791
rect 1984 6771 2604 6781
rect 2614 6771 2634 6781
rect 2654 6771 2854 6781
rect 1994 6761 2874 6771
rect 1994 6751 2894 6761
rect 1994 6741 2944 6751
rect 1994 6731 2954 6741
rect 1994 6721 2964 6731
rect 1974 6711 2974 6721
rect 1964 6701 2644 6711
rect 2674 6701 2974 6711
rect 1954 6691 2614 6701
rect 2684 6691 2924 6701
rect 1944 6671 2614 6691
rect 2754 6681 2924 6691
rect 2774 6671 2904 6681
rect 1934 6661 2624 6671
rect 2794 6661 2904 6671
rect 1924 6651 2634 6661
rect 2834 6651 2904 6661
rect 1914 6641 2634 6651
rect 2854 6641 2914 6651
rect 3714 6641 3734 6651
rect 1894 6621 2564 6641
rect 2574 6631 2634 6641
rect 2884 6631 2934 6641
rect 3714 6631 3764 6641
rect 2584 6621 2634 6631
rect 2894 6621 2934 6631
rect 3724 6621 3764 6631
rect 1894 6611 2554 6621
rect 2614 6611 2634 6621
rect 2914 6611 2934 6621
rect 3714 6611 3814 6621
rect 1874 6591 2544 6611
rect 3674 6601 3814 6611
rect 3674 6591 3854 6601
rect 1894 6581 2224 6591
rect 2264 6581 2554 6591
rect 3694 6581 3874 6591
rect 1894 6571 2214 6581
rect 1864 6561 2204 6571
rect 2274 6561 2554 6581
rect 3014 6571 3064 6581
rect 3704 6571 3884 6581
rect 3014 6561 3074 6571
rect 3724 6561 3884 6571
rect 1864 6551 2134 6561
rect 2144 6551 2204 6561
rect 1864 6531 2204 6551
rect 1854 6521 2204 6531
rect 2244 6521 2254 6531
rect 1774 6511 1784 6521
rect 1844 6511 2204 6521
rect 2234 6511 2254 6521
rect 2284 6521 2554 6561
rect 3024 6551 3084 6561
rect 3284 6551 3324 6561
rect 3724 6551 3914 6561
rect 3054 6541 3094 6551
rect 3064 6531 3104 6541
rect 3284 6531 3344 6551
rect 3404 6541 3414 6551
rect 3444 6541 3464 6551
rect 3734 6541 3924 6551
rect 3434 6531 3484 6541
rect 3754 6531 3934 6541
rect 3084 6521 3094 6531
rect 2284 6511 2564 6521
rect 3294 6511 3334 6531
rect 3424 6521 3494 6531
rect 3754 6521 3974 6531
rect 3424 6511 3514 6521
rect 3784 6511 3974 6521
rect 1764 6501 1794 6511
rect 1844 6501 2202 6511
rect 2244 6501 2254 6511
rect 1754 6491 1804 6501
rect 1844 6491 2184 6501
rect 2294 6491 2574 6511
rect 3294 6501 3344 6511
rect 3424 6501 3454 6511
rect 3464 6501 3534 6511
rect 3794 6501 3984 6511
rect 3304 6491 3354 6501
rect 3474 6491 3554 6501
rect 3814 6491 4014 6501
rect 1754 6481 1814 6491
rect 1834 6481 2194 6491
rect 2294 6481 2584 6491
rect 3324 6481 3364 6491
rect 3484 6481 3564 6491
rect 3824 6481 4034 6491
rect 1754 6471 2194 6481
rect 2284 6471 2404 6481
rect 2434 6471 2604 6481
rect 3334 6471 3374 6481
rect 3504 6471 3584 6481
rect 3834 6471 4044 6481
rect 1744 6461 2194 6471
rect 2294 6461 2394 6471
rect 2434 6461 2614 6471
rect 1744 6451 2074 6461
rect 1734 6441 2034 6451
rect 2054 6441 2074 6451
rect 1724 6431 1984 6441
rect 2004 6431 2034 6441
rect 1714 6421 1984 6431
rect 2014 6421 2034 6431
rect 2064 6421 2074 6441
rect 2094 6431 2184 6461
rect 2294 6451 2384 6461
rect 2424 6451 2614 6461
rect 3354 6461 3374 6471
rect 3514 6461 3594 6471
rect 3844 6461 4064 6471
rect 3354 6451 3384 6461
rect 3524 6451 3594 6461
rect 3854 6451 4084 6461
rect 2304 6441 2374 6451
rect 2414 6441 2594 6451
rect 3374 6441 3414 6451
rect 3524 6441 3574 6451
rect 3864 6441 4114 6451
rect 2274 6431 2284 6441
rect 2304 6431 2364 6441
rect 2404 6431 2474 6441
rect 2104 6421 2184 6431
rect 2264 6421 2284 6431
rect 2294 6421 2354 6431
rect 2394 6421 2464 6431
rect 1704 6411 1984 6421
rect 2104 6411 2174 6421
rect 2294 6411 2344 6421
rect 1694 6391 1984 6411
rect 1684 6381 1714 6391
rect 1724 6381 1984 6391
rect 2114 6381 2174 6411
rect 2284 6401 2344 6411
rect 2384 6411 2444 6421
rect 2484 6411 2564 6441
rect 3384 6431 3424 6441
rect 3534 6431 3564 6441
rect 3874 6431 4134 6441
rect 3394 6421 3434 6431
rect 3554 6421 3604 6431
rect 3874 6421 4154 6431
rect 3404 6411 3444 6421
rect 2384 6401 2424 6411
rect 2474 6401 2574 6411
rect 3414 6401 3454 6411
rect 3564 6401 3614 6421
rect 3874 6411 4174 6421
rect 3624 6401 3634 6411
rect 3914 6401 4174 6411
rect 2284 6391 2334 6401
rect 2354 6391 2364 6401
rect 2394 6391 2404 6401
rect 2274 6381 2324 6391
rect 1684 6371 1704 6381
rect 1734 6371 1974 6381
rect 1664 6351 1674 6361
rect 1744 6351 1964 6371
rect 2114 6361 2164 6381
rect 2264 6371 2314 6381
rect 1654 6331 1674 6351
rect 1754 6341 1954 6351
rect 1764 6331 1954 6341
rect 2114 6331 2154 6361
rect 2264 6351 2324 6371
rect 2354 6361 2374 6391
rect 2464 6381 2574 6401
rect 3424 6391 3474 6401
rect 3574 6391 3584 6401
rect 3424 6381 3494 6391
rect 3594 6381 3644 6401
rect 3904 6391 4204 6401
rect 3924 6381 4214 6391
rect 2464 6371 2584 6381
rect 2454 6361 2594 6371
rect 2704 6361 2734 6381
rect 3434 6371 3504 6381
rect 3594 6371 3664 6381
rect 3934 6371 4224 6381
rect 3434 6361 3524 6371
rect 3624 6361 3664 6371
rect 3944 6361 4224 6371
rect 2454 6351 2604 6361
rect 2704 6351 2744 6361
rect 3444 6351 3524 6361
rect 3634 6351 3664 6361
rect 3954 6351 4234 6361
rect 2274 6341 2324 6351
rect 2464 6341 2614 6351
rect 2274 6331 2314 6341
rect 2454 6331 2614 6341
rect 2724 6341 2754 6351
rect 3284 6341 3304 6351
rect 3454 6341 3534 6351
rect 3724 6341 3754 6351
rect 3964 6341 4244 6351
rect 2724 6331 2774 6341
rect 3284 6331 3324 6341
rect 3474 6331 3544 6341
rect 3724 6331 3774 6341
rect 3974 6331 4244 6341
rect 1644 6321 1674 6331
rect 1774 6321 1944 6331
rect 2124 6321 2144 6331
rect 2244 6321 2304 6331
rect 2444 6321 2614 6331
rect 2734 6321 2784 6331
rect 3164 6321 3204 6331
rect 3284 6321 3344 6331
rect 1644 6311 1664 6321
rect 1774 6311 1814 6321
rect 1824 6311 1934 6321
rect 2224 6311 2284 6321
rect 2434 6311 2625 6321
rect 2774 6311 2844 6321
rect 2864 6311 2894 6321
rect 2964 6311 2984 6321
rect 3164 6311 3214 6321
rect 3264 6311 3344 6321
rect 3484 6321 3594 6331
rect 3724 6321 3824 6331
rect 3984 6321 4254 6331
rect 3484 6311 3604 6321
rect 3724 6311 3834 6321
rect 4014 6311 4254 6321
rect 1704 6301 1724 6311
rect 1774 6301 1804 6311
rect 1824 6301 1924 6311
rect 2224 6301 2274 6311
rect 2424 6301 2654 6311
rect 2784 6301 2904 6311
rect 2964 6301 3014 6311
rect 3174 6301 3364 6311
rect 3494 6301 3614 6311
rect 3734 6301 3844 6311
rect 4024 6301 4284 6311
rect 1704 6281 1734 6301
rect 1714 6271 1734 6281
rect 1824 6291 1914 6301
rect 2224 6291 2244 6301
rect 2264 6291 2274 6301
rect 2414 6291 2654 6301
rect 2794 6291 2914 6301
rect 2974 6291 3024 6301
rect 3174 6291 3204 6301
rect 3214 6291 3374 6301
rect 3504 6291 3634 6301
rect 3744 6291 3854 6301
rect 4024 6291 4334 6301
rect 1824 6271 1904 6291
rect 2414 6281 2664 6291
rect 2804 6281 2924 6291
rect 2974 6281 3034 6291
rect 3174 6281 3394 6291
rect 3514 6281 3644 6291
rect 3754 6281 3864 6291
rect 4034 6281 4344 6291
rect 2214 6271 2224 6281
rect 2414 6271 2524 6281
rect 1814 6251 1904 6271
rect 1634 6231 1654 6241
rect 1724 6231 1734 6241
rect 1634 6201 1664 6231
rect 1714 6221 1734 6231
rect 1804 6231 1894 6251
rect 2194 6241 2224 6271
rect 2304 6251 2314 6271
rect 2404 6261 2514 6271
rect 2394 6241 2514 6261
rect 2534 6251 2674 6281
rect 2814 6271 2924 6281
rect 2984 6271 3054 6281
rect 3174 6271 3414 6281
rect 3534 6271 3664 6281
rect 3764 6271 3884 6281
rect 2834 6261 2934 6271
rect 2994 6261 3054 6271
rect 3194 6261 3204 6271
rect 3214 6261 3424 6271
rect 3544 6261 3674 6271
rect 3784 6261 3894 6271
rect 4044 6261 4304 6281
rect 4324 6271 4364 6281
rect 4334 6261 4374 6271
rect 2844 6251 2944 6261
rect 3004 6251 3084 6261
rect 3194 6251 3444 6261
rect 3554 6251 3684 6261
rect 3794 6251 3904 6261
rect 4054 6251 4364 6261
rect 2194 6231 2214 6241
rect 2384 6231 2514 6241
rect 1804 6211 1884 6231
rect 2384 6221 2504 6231
rect 2374 6211 2394 6221
rect 1804 6201 1874 6211
rect 2364 6201 2394 6211
rect 1644 6181 1674 6201
rect 1804 6191 1864 6201
rect 1714 6181 1724 6191
rect 1794 6181 1854 6191
rect 2164 6181 2174 6201
rect 2364 6181 2384 6201
rect 2414 6181 2504 6221
rect 2524 6221 2704 6251
rect 2864 6241 2954 6251
rect 3014 6241 3104 6251
rect 2874 6231 2954 6241
rect 3024 6231 3104 6241
rect 3184 6241 3454 6251
rect 3554 6241 3694 6251
rect 3794 6241 3914 6251
rect 4074 6241 4374 6251
rect 3184 6231 3464 6241
rect 3554 6231 3714 6241
rect 3804 6231 3924 6241
rect 4014 6231 4024 6241
rect 4094 6231 4374 6241
rect 2884 6221 2964 6231
rect 3034 6221 3124 6231
rect 3144 6221 3154 6231
rect 3174 6221 3474 6231
rect 3564 6221 3734 6231
rect 3814 6221 3974 6231
rect 3984 6221 4034 6231
rect 4134 6221 4384 6231
rect 2524 6211 2714 6221
rect 2894 6211 2964 6221
rect 3064 6211 3494 6221
rect 3574 6211 3734 6221
rect 3824 6211 4034 6221
rect 4144 6211 4394 6221
rect 2524 6201 2724 6211
rect 2904 6201 2954 6211
rect 3074 6201 3514 6211
rect 3584 6201 3754 6211
rect 3834 6201 4044 6211
rect 4134 6201 4394 6211
rect 2524 6181 2684 6201
rect 2704 6191 2724 6201
rect 3094 6191 3514 6201
rect 3594 6191 3764 6201
rect 3844 6191 4054 6201
rect 4124 6191 4384 6201
rect 1634 6171 1724 6181
rect 1624 6161 1714 6171
rect 1784 6161 1844 6181
rect 2364 6171 2374 6181
rect 2404 6161 2494 6181
rect 1624 6151 1704 6161
rect 1634 6141 1704 6151
rect 1784 6141 1834 6161
rect 2194 6151 2204 6161
rect 2394 6151 2494 6161
rect 2174 6141 2184 6151
rect 2194 6141 2214 6151
rect 1624 6131 1714 6141
rect 1764 6131 1824 6141
rect 2164 6131 2184 6141
rect 1624 6111 1724 6131
rect 1754 6121 1814 6131
rect 1744 6111 1784 6121
rect 2334 6111 2354 6141
rect 1624 6101 1774 6111
rect 2324 6101 2354 6111
rect 2384 6131 2424 6151
rect 2454 6141 2494 6151
rect 2524 6171 2694 6181
rect 2704 6171 2734 6191
rect 3094 6181 3234 6191
rect 3264 6181 3524 6191
rect 3604 6181 3764 6191
rect 3854 6181 4074 6191
rect 4134 6181 4154 6191
rect 4174 6181 4384 6191
rect 3104 6171 3244 6181
rect 3274 6171 3524 6181
rect 3624 6171 3784 6181
rect 3864 6171 3894 6181
rect 3954 6171 4074 6181
rect 2524 6161 2744 6171
rect 3094 6161 3124 6171
rect 3134 6161 3254 6171
rect 3284 6161 3524 6171
rect 3634 6161 3794 6171
rect 3904 6161 3924 6171
rect 3944 6161 4104 6171
rect 4224 6161 4384 6181
rect 2524 6151 2754 6161
rect 3094 6151 3114 6161
rect 3154 6151 3264 6161
rect 3294 6151 3534 6161
rect 3654 6151 3804 6161
rect 3884 6151 4124 6161
rect 4234 6151 4394 6161
rect 2524 6141 2574 6151
rect 2604 6141 2764 6151
rect 3096 6150 3274 6151
rect 2454 6131 2484 6141
rect 2524 6131 2564 6141
rect 2384 6111 2414 6131
rect 2454 6121 2474 6131
rect 2444 6111 2474 6121
rect 2524 6111 2544 6131
rect 2594 6121 2764 6141
rect 3104 6141 3274 6150
rect 3304 6141 3534 6151
rect 3674 6141 3814 6151
rect 3884 6141 4144 6151
rect 4244 6141 4424 6151
rect 3104 6131 3284 6141
rect 3314 6131 3554 6141
rect 3684 6131 3854 6141
rect 3884 6131 4154 6141
rect 4264 6131 4424 6141
rect 2584 6120 2764 6121
rect 2574 6111 2764 6120
rect 3094 6121 3294 6131
rect 3334 6121 3584 6131
rect 3684 6121 3864 6131
rect 3894 6121 4154 6131
rect 4294 6121 4424 6131
rect 3094 6111 3304 6121
rect 3354 6111 3594 6121
rect 3694 6111 3874 6121
rect 3904 6111 4174 6121
rect 4294 6111 4434 6121
rect 2384 6101 2404 6111
rect 2434 6101 2464 6111
rect 2554 6108 2774 6111
rect 2554 6101 2584 6108
rect 2604 6101 2774 6108
rect 3104 6101 3344 6111
rect 1614 6091 1734 6101
rect 1604 6081 1734 6091
rect 1594 6071 1724 6081
rect 1584 6061 1724 6071
rect 1584 6021 1764 6061
rect 2314 6051 2344 6101
rect 2374 6091 2394 6101
rect 2434 6091 2454 6101
rect 2554 6091 2574 6101
rect 2604 6091 2784 6101
rect 3114 6091 3344 6101
rect 3364 6091 3594 6111
rect 3714 6101 3894 6111
rect 3904 6102 4194 6111
rect 3904 6101 4206 6102
rect 3724 6091 4206 6101
rect 4294 6101 4444 6111
rect 4294 6091 4344 6101
rect 4384 6091 4454 6101
rect 2364 6071 2394 6091
rect 2544 6071 2564 6091
rect 2314 6031 2334 6051
rect 2364 6041 2384 6071
rect 2554 6061 2564 6071
rect 2614 6081 2794 6091
rect 3124 6081 3354 6091
rect 3364 6081 3624 6091
rect 3734 6081 4174 6091
rect 4185 6090 4214 6091
rect 4194 6081 4214 6090
rect 4304 6081 4354 6091
rect 4394 6081 4464 6091
rect 2614 6071 2804 6081
rect 3134 6071 3634 6081
rect 3744 6071 4164 6081
rect 4194 6071 4204 6081
rect 2614 6061 2824 6071
rect 3144 6061 3644 6071
rect 2624 6051 2834 6061
rect 3154 6051 3644 6061
rect 3754 6061 4204 6071
rect 3754 6051 4224 6061
rect 2364 6031 2374 6041
rect 2554 6031 2564 6051
rect 2654 6041 2834 6051
rect 3184 6041 3644 6051
rect 3734 6041 3764 6051
rect 2664 6031 2734 6041
rect 2744 6031 2874 6041
rect 3194 6031 3684 6041
rect 1574 6001 1764 6021
rect 2354 6011 2374 6031
rect 2344 6001 2374 6011
rect 2684 6021 2734 6031
rect 2754 6021 2884 6031
rect 3214 6021 3694 6031
rect 3724 6021 3764 6041
rect 3794 6041 3814 6051
rect 3824 6041 4254 6051
rect 4324 6041 4374 6081
rect 4404 6071 4464 6081
rect 4414 6061 4464 6071
rect 4414 6051 4474 6061
rect 4424 6041 4474 6051
rect 3794 6021 3804 6041
rect 3834 6031 4264 6041
rect 4334 6031 4374 6041
rect 4434 6031 4474 6041
rect 3834 6021 3864 6031
rect 3934 6021 4274 6031
rect 4364 6021 4384 6031
rect 2684 6001 2744 6021
rect 2754 6011 2894 6021
rect 3224 6011 3764 6021
rect 3934 6011 4284 6021
rect 4364 6011 4394 6021
rect 2763 6001 2924 6011
rect 3234 6001 3774 6011
rect 3934 6001 4184 6011
rect 4244 6001 4314 6011
rect 4454 6001 4484 6031
rect 1574 5991 1754 6001
rect 2354 5991 2364 6001
rect 2694 5991 2754 6001
rect 2763 5991 2954 6001
rect 3244 5991 3784 6001
rect 3944 5991 3974 6001
rect 3984 5991 4164 6001
rect 4264 5991 4324 6001
rect 1574 5981 1744 5991
rect 2654 5981 2664 5991
rect 2694 5981 2774 5991
rect 2794 5981 2974 5991
rect 3264 5981 3804 5991
rect 3954 5981 4144 5991
rect 4274 5981 4324 5991
rect 1574 5971 1614 5981
rect 1624 5971 1744 5981
rect 1574 5951 1744 5971
rect 2694 5971 2994 5981
rect 3274 5971 3834 5981
rect 3974 5971 4124 5981
rect 4304 5971 4324 5981
rect 2694 5961 3004 5971
rect 3284 5961 3844 5971
rect 3984 5961 4154 5971
rect 2684 5951 3014 5961
rect 3284 5951 3854 5961
rect 3994 5951 4164 5961
rect 4374 5951 4394 5961
rect 1584 5941 1734 5951
rect 1604 5921 1734 5941
rect 1764 5941 1784 5951
rect 2684 5941 2804 5951
rect 2814 5941 3034 5951
rect 3304 5941 3864 5951
rect 4004 5941 4164 5951
rect 4354 5941 4424 5951
rect 1764 5931 1774 5941
rect 2694 5931 3054 5941
rect 3324 5931 3904 5941
rect 4024 5931 4164 5941
rect 4364 5931 4454 5941
rect 2704 5921 3064 5931
rect 3144 5921 3164 5931
rect 3334 5921 3904 5931
rect 4064 5921 4174 5931
rect 4374 5921 4464 5931
rect 1614 5901 1744 5921
rect 2174 5901 2194 5921
rect 1614 5891 1734 5901
rect 2174 5891 2184 5901
rect 1624 5881 1694 5891
rect 1614 5871 1684 5881
rect 2164 5871 2174 5881
rect 2454 5871 2464 5921
rect 2704 5911 3094 5921
rect 3134 5911 3204 5921
rect 3334 5911 3934 5921
rect 4094 5911 4214 5921
rect 2704 5901 2844 5911
rect 2854 5901 3214 5911
rect 3334 5910 3954 5911
rect 3334 5901 3464 5910
rect 3494 5901 3954 5910
rect 4104 5901 4224 5911
rect 2704 5891 2834 5901
rect 2854 5891 3224 5901
rect 3344 5891 3474 5901
rect 3504 5891 3974 5901
rect 4124 5891 4224 5901
rect 4384 5891 4464 5921
rect 2704 5871 3254 5891
rect 3374 5881 3484 5891
rect 3514 5881 3994 5891
rect 4134 5881 4224 5891
rect 3384 5871 3494 5881
rect 3524 5871 4004 5881
rect 4144 5871 4224 5881
rect 4284 5871 4304 5881
rect 4394 5871 4464 5891
rect 1614 5861 1674 5871
rect 2074 5861 2084 5871
rect 2154 5861 2184 5871
rect 1624 5841 1664 5861
rect 2064 5851 2084 5861
rect 2144 5851 2184 5861
rect 2454 5851 2474 5871
rect 2704 5861 2774 5871
rect 2784 5861 3264 5871
rect 3394 5861 3504 5871
rect 3534 5861 4004 5871
rect 4184 5861 4204 5871
rect 2704 5851 3284 5861
rect 3404 5851 3514 5861
rect 2054 5841 2094 5851
rect 1634 5831 1664 5841
rect 1624 5821 1664 5831
rect 2044 5821 2094 5841
rect 2144 5831 2174 5851
rect 2464 5841 2484 5851
rect 2704 5841 3294 5851
rect 3404 5841 3524 5851
rect 3544 5841 4004 5861
rect 4264 5851 4314 5871
rect 4404 5861 4464 5871
rect 4414 5851 4464 5861
rect 4414 5841 4454 5851
rect 2134 5821 2174 5831
rect 1624 5811 1654 5821
rect 2044 5811 2084 5821
rect 1624 5801 1644 5811
rect 2044 5801 2064 5811
rect 1614 5781 1654 5801
rect 2034 5781 2074 5801
rect 1614 5771 1664 5781
rect 1614 5751 1654 5771
rect 1774 5761 1784 5771
rect 1764 5751 1784 5761
rect 1614 5741 1644 5751
rect 1624 5731 1644 5741
rect 1634 5711 1644 5731
rect 1754 5721 1784 5751
rect 2044 5761 2074 5781
rect 2044 5731 2084 5761
rect 1764 5711 1784 5721
rect 2054 5711 2084 5731
rect 1754 5701 1784 5711
rect 1634 5681 1654 5691
rect 1744 5681 1784 5701
rect 2064 5701 2084 5711
rect 2144 5701 2174 5821
rect 2454 5821 2494 5841
rect 2534 5831 2554 5841
rect 2704 5831 3314 5841
rect 3414 5831 3534 5841
rect 3574 5831 4004 5841
rect 4284 5831 4334 5841
rect 2454 5811 2504 5821
rect 2534 5811 2564 5831
rect 2714 5821 3324 5831
rect 3424 5821 3544 5831
rect 3584 5821 4014 5831
rect 4284 5821 4324 5831
rect 2714 5811 3344 5821
rect 3434 5811 3544 5821
rect 3594 5811 4024 5821
rect 2464 5791 2504 5811
rect 2544 5801 2554 5811
rect 2724 5801 3344 5811
rect 3444 5801 3564 5811
rect 2544 5791 2604 5801
rect 2464 5781 2514 5791
rect 2554 5781 2604 5791
rect 2734 5791 3364 5801
rect 3464 5791 3564 5801
rect 3604 5801 4044 5811
rect 3604 5791 4074 5801
rect 2734 5781 3374 5791
rect 2464 5771 2524 5781
rect 2554 5771 2614 5781
rect 2744 5771 3274 5781
rect 3294 5771 3374 5781
rect 3484 5781 3564 5791
rect 3614 5781 4074 5791
rect 3484 5771 3574 5781
rect 3624 5771 4084 5781
rect 2474 5761 2524 5771
rect 2564 5761 2624 5771
rect 2744 5761 3394 5771
rect 3484 5761 3584 5771
rect 3624 5761 4104 5771
rect 2334 5731 2354 5751
rect 2484 5741 2534 5761
rect 2574 5751 2634 5761
rect 2564 5741 2634 5751
rect 2754 5751 3294 5761
rect 3314 5751 3414 5761
rect 3514 5751 3614 5761
rect 3634 5751 4114 5761
rect 2754 5741 3304 5751
rect 3324 5741 3424 5751
rect 3524 5741 4114 5751
rect 2494 5721 2544 5741
rect 2574 5721 2644 5741
rect 2754 5721 3354 5741
rect 3384 5731 3424 5741
rect 3534 5731 4134 5741
rect 3414 5721 3424 5731
rect 3544 5721 3654 5731
rect 3674 5721 4144 5731
rect 2364 5701 2394 5721
rect 2494 5711 2554 5721
rect 2064 5681 2094 5701
rect 2144 5691 2194 5701
rect 2364 5691 2414 5701
rect 2504 5691 2564 5711
rect 1624 5651 1664 5681
rect 1744 5661 1774 5681
rect 2064 5661 2104 5681
rect 2144 5671 2204 5691
rect 2384 5681 2414 5691
rect 2514 5681 2564 5691
rect 2594 5701 2664 5721
rect 2754 5711 3364 5721
rect 2754 5701 3374 5711
rect 2594 5681 2674 5701
rect 2754 5691 3404 5701
rect 3434 5691 3464 5721
rect 3554 5711 3644 5721
rect 3684 5711 4154 5721
rect 3554 5701 3654 5711
rect 3674 5701 4144 5711
rect 4404 5701 4424 5711
rect 3554 5691 4144 5701
rect 4394 5691 4444 5701
rect 2764 5681 3484 5691
rect 3564 5681 4154 5691
rect 4404 5681 4454 5691
rect 2384 5671 2424 5681
rect 2514 5671 2574 5681
rect 2604 5671 2684 5681
rect 2774 5671 3504 5681
rect 3574 5671 4154 5681
rect 4324 5671 4334 5681
rect 4394 5671 4454 5681
rect 2154 5661 2194 5671
rect 2394 5661 2454 5671
rect 2514 5661 2584 5671
rect 2624 5661 2684 5671
rect 2784 5661 3534 5671
rect 3584 5661 4164 5671
rect 4304 5661 4354 5671
rect 4394 5661 4444 5671
rect 1744 5651 1764 5661
rect 1624 5641 1674 5651
rect 1714 5641 1764 5651
rect 1624 5631 1684 5641
rect 1704 5631 1764 5641
rect 1624 5621 1764 5631
rect 1614 5611 1764 5621
rect 1944 5641 1974 5651
rect 2064 5641 2114 5661
rect 1944 5621 1984 5641
rect 2074 5621 2114 5641
rect 1944 5611 2024 5621
rect 1614 5601 1744 5611
rect 1944 5601 2034 5611
rect 2064 5601 2114 5621
rect 2164 5651 2204 5661
rect 2404 5651 2474 5661
rect 2524 5651 2594 5661
rect 2624 5651 2704 5661
rect 2794 5651 3094 5661
rect 3104 5651 3544 5661
rect 3594 5651 4094 5661
rect 4114 5651 4174 5661
rect 4304 5651 4364 5661
rect 4404 5651 4444 5661
rect 2164 5641 2214 5651
rect 2404 5641 2484 5651
rect 2534 5641 2604 5651
rect 2634 5641 2714 5651
rect 2804 5641 3094 5651
rect 3114 5641 3554 5651
rect 3594 5641 4104 5651
rect 4124 5643 4194 5651
rect 4124 5641 4143 5643
rect 4155 5641 4194 5643
rect 4304 5641 4384 5651
rect 4394 5641 4444 5651
rect 2164 5611 2224 5641
rect 2404 5631 2494 5641
rect 2534 5631 2614 5641
rect 2644 5631 2724 5641
rect 2804 5631 3104 5641
rect 3124 5631 3564 5641
rect 3604 5631 4104 5641
rect 2414 5621 2504 5631
rect 2534 5621 2624 5631
rect 2634 5621 2734 5631
rect 2814 5621 3114 5631
rect 3134 5621 3154 5631
rect 3164 5621 3574 5631
rect 3594 5621 4124 5631
rect 4134 5621 4143 5631
rect 4155 5622 4204 5641
rect 4161 5621 4204 5622
rect 4314 5631 4444 5641
rect 4314 5621 4434 5631
rect 2424 5611 2514 5621
rect 2554 5611 2744 5621
rect 2824 5611 3124 5621
rect 3174 5619 4143 5621
rect 3174 5611 4144 5619
rect 4164 5611 4204 5621
rect 4334 5611 4434 5621
rect 2164 5601 2234 5611
rect 1614 5581 1754 5601
rect 1944 5581 2044 5601
rect 1604 5571 1744 5581
rect 1614 5551 1734 5571
rect 1944 5561 2054 5581
rect 2074 5571 2114 5601
rect 2174 5591 2234 5601
rect 2184 5581 2234 5591
rect 2254 5601 2274 5611
rect 2434 5601 2524 5611
rect 2544 5601 2644 5611
rect 2654 5601 2764 5611
rect 2844 5601 3134 5611
rect 3174 5601 4154 5611
rect 4194 5601 4214 5611
rect 4344 5601 4434 5611
rect 2254 5591 2284 5601
rect 2434 5591 2534 5601
rect 2554 5591 2644 5601
rect 2664 5591 2774 5601
rect 2844 5591 3144 5601
rect 3164 5591 4174 5601
rect 4194 5591 4224 5601
rect 4334 5591 4434 5601
rect 2254 5581 2294 5591
rect 2444 5581 2654 5591
rect 2084 5561 2124 5571
rect 2184 5561 2224 5581
rect 2264 5571 2314 5581
rect 2464 5571 2654 5581
rect 2674 5581 2784 5591
rect 2844 5581 2854 5591
rect 2864 5581 3174 5591
rect 3184 5581 4174 5591
rect 4314 5581 4354 5591
rect 4384 5581 4434 5591
rect 2674 5571 2754 5581
rect 2764 5571 2804 5581
rect 2844 5571 4184 5581
rect 4304 5571 4424 5581
rect 2264 5561 2334 5571
rect 2474 5561 2664 5571
rect 2674 5561 2814 5571
rect 2854 5561 4194 5571
rect 4314 5561 4424 5571
rect 1774 5551 1784 5561
rect 1944 5551 2064 5561
rect 2084 5551 2134 5561
rect 2194 5551 2234 5561
rect 2264 5551 2344 5561
rect 2494 5551 2814 5561
rect 2844 5551 3204 5561
rect 1604 5541 1734 5551
rect 1754 5541 1784 5551
rect 1894 5541 1904 5551
rect 1944 5541 2074 5551
rect 2084 5541 2144 5551
rect 1604 5521 1784 5541
rect 1944 5531 2144 5541
rect 2194 5531 2254 5551
rect 2284 5541 2354 5551
rect 2504 5541 2694 5551
rect 2704 5541 3204 5551
rect 3214 5551 4204 5561
rect 4304 5551 4424 5561
rect 3214 5541 4214 5551
rect 4304 5541 4414 5551
rect 2284 5531 2374 5541
rect 2534 5531 2854 5541
rect 2864 5531 3204 5541
rect 3224 5531 4224 5541
rect 1934 5521 2154 5531
rect 2204 5521 2264 5531
rect 2294 5521 2394 5531
rect 2554 5521 3214 5531
rect 1604 5491 1794 5521
rect 1934 5511 2164 5521
rect 2214 5511 2264 5521
rect 2304 5511 2414 5521
rect 2624 5511 3214 5521
rect 3234 5521 4244 5531
rect 3234 5511 4254 5521
rect 4314 5511 4414 5541
rect 1964 5501 2174 5511
rect 2214 5501 2274 5511
rect 2314 5501 2424 5511
rect 2634 5501 3224 5511
rect 3234 5501 4274 5511
rect 1604 5471 1804 5491
rect 1924 5481 2204 5501
rect 2224 5491 2294 5501
rect 2244 5481 2294 5491
rect 1914 5471 2204 5481
rect 1604 5451 1814 5471
rect 1604 5411 1824 5451
rect 1924 5441 2204 5471
rect 2214 5471 2234 5481
rect 2254 5471 2294 5481
rect 2324 5491 2484 5501
rect 2634 5491 4284 5501
rect 4324 5491 4414 5511
rect 2324 5481 2494 5491
rect 2624 5481 4294 5491
rect 2324 5471 2554 5481
rect 2564 5471 3794 5481
rect 3804 5471 4314 5481
rect 4334 5471 4414 5491
rect 2214 5451 2244 5471
rect 2264 5461 2284 5471
rect 2324 5461 2764 5471
rect 2344 5460 2774 5461
rect 2784 5460 4414 5471
rect 2344 5451 4414 5460
rect 2214 5441 2254 5451
rect 2284 5441 2294 5451
rect 2354 5441 2784 5451
rect 1924 5431 2304 5441
rect 2364 5431 2794 5441
rect 2824 5431 4414 5451
rect 1924 5421 2314 5431
rect 2324 5421 2344 5431
rect 2364 5421 2804 5431
rect 2814 5421 4414 5431
rect 1924 5411 2344 5421
rect 1604 5401 1834 5411
rect 1924 5401 2354 5411
rect 2414 5401 4414 5421
rect 1614 5381 1834 5401
rect 1934 5391 2364 5401
rect 2414 5391 2834 5401
rect 2854 5391 4414 5401
rect 1934 5381 2374 5391
rect 2414 5381 2444 5391
rect 1614 5371 1844 5381
rect 1944 5371 2434 5381
rect 2464 5371 4414 5391
rect 1624 5341 1854 5371
rect 1944 5361 4414 5371
rect 1954 5351 4414 5361
rect 1954 5341 4424 5351
rect 1624 5321 1864 5341
rect 1964 5321 4424 5341
rect 1624 5301 1874 5321
rect 1974 5311 4424 5321
rect 1984 5301 4434 5311
rect 1624 5281 1884 5301
rect 1994 5291 2544 5301
rect 1994 5281 2534 5291
rect 2554 5281 4434 5301
rect 1624 5261 1894 5281
rect 2014 5271 2223 5281
rect 2234 5271 4434 5281
rect 4594 5271 4614 5281
rect 1944 5261 1954 5271
rect 2004 5261 2204 5271
rect 2214 5261 2224 5271
rect 2244 5261 2274 5271
rect 2284 5261 4424 5271
rect 4594 5261 4634 5271
rect 1624 5241 1904 5261
rect 1934 5251 1974 5261
rect 2004 5251 2224 5261
rect 2254 5251 2264 5261
rect 2314 5251 2384 5261
rect 2404 5251 4414 5261
rect 4574 5251 4634 5261
rect 1944 5241 1974 5251
rect 1984 5241 2124 5251
rect 2154 5241 2234 5251
rect 2344 5241 2374 5251
rect 2444 5241 4404 5251
rect 4574 5241 4624 5251
rect 1624 5221 1934 5241
rect 1944 5231 2114 5241
rect 2154 5231 2184 5241
rect 2214 5231 2234 5241
rect 2464 5231 4404 5241
rect 4584 5231 4594 5241
rect 4604 5231 4624 5241
rect 1944 5221 2134 5231
rect 2544 5221 4384 5231
rect 1624 5191 2154 5221
rect 2554 5211 4384 5221
rect 2564 5201 2594 5211
rect 2624 5201 4374 5211
rect 2624 5191 4364 5201
rect 1624 5181 2094 5191
rect 2124 5181 2144 5191
rect 2614 5181 4364 5191
rect 1624 5171 2104 5181
rect 2614 5171 2634 5181
rect 2644 5171 4364 5181
rect 1624 5161 2114 5171
rect 2604 5161 2624 5171
rect 2654 5161 2804 5171
rect 1624 5151 2144 5161
rect 2604 5151 2634 5161
rect 1634 5141 2154 5151
rect 2624 5141 2634 5151
rect 2644 5151 2804 5161
rect 2814 5151 4354 5171
rect 2644 5141 2764 5151
rect 2824 5141 4344 5151
rect 1634 5131 2164 5141
rect 2654 5131 2764 5141
rect 1644 5121 2174 5131
rect 1644 5111 2054 5121
rect 2074 5111 2154 5121
rect 1584 5081 1614 5111
rect 1644 5101 2044 5111
rect 2084 5101 2114 5111
rect 2164 5101 2194 5111
rect 2364 5101 2384 5131
rect 2684 5121 2764 5131
rect 2704 5111 2734 5121
rect 2754 5101 2764 5121
rect 2814 5111 2854 5141
rect 2864 5131 4344 5141
rect 2874 5121 4314 5131
rect 2874 5111 4284 5121
rect 2874 5101 4134 5111
rect 4144 5101 4284 5111
rect 1654 5091 2044 5101
rect 2174 5091 2184 5101
rect 2894 5091 4134 5101
rect 4154 5091 4284 5101
rect 1664 5081 2024 5091
rect 2914 5081 4144 5091
rect 1584 5051 1624 5081
rect 1674 5071 2014 5081
rect 2934 5071 4144 5081
rect 4164 5081 4274 5091
rect 4164 5071 4264 5081
rect 1674 5051 2004 5071
rect 2374 5061 2404 5071
rect 2954 5061 4154 5071
rect 4164 5061 4254 5071
rect 1574 5021 1624 5051
rect 1684 5041 2004 5051
rect 2324 5051 2464 5061
rect 2504 5051 2524 5061
rect 2974 5051 4254 5061
rect 2324 5041 2584 5051
rect 2984 5041 4184 5051
rect 1684 5031 1994 5041
rect 2314 5031 2644 5041
rect 3024 5031 4184 5041
rect 4194 5041 4244 5051
rect 4194 5031 4234 5041
rect 1564 4991 1624 5021
rect 1704 5021 1984 5031
rect 2224 5021 2234 5031
rect 2314 5021 2664 5031
rect 3104 5021 4224 5031
rect 1704 5011 1974 5021
rect 2214 5011 2274 5021
rect 2354 5011 2684 5021
rect 3174 5011 3194 5021
rect 3204 5011 4204 5021
rect 1554 4981 1624 4991
rect 1694 5001 1974 5011
rect 2234 5001 2264 5011
rect 2394 5001 2704 5011
rect 2714 5001 2734 5011
rect 3214 5001 4194 5011
rect 1694 4991 1964 5001
rect 2404 4991 2754 5001
rect 3224 4991 4184 5001
rect 1694 4981 1954 4991
rect 2434 4981 2464 4991
rect 2504 4981 2764 4991
rect 3234 4981 4154 4991
rect 1544 4971 1624 4981
rect 1704 4971 1954 4981
rect 2534 4971 2774 4981
rect 3254 4971 4124 4981
rect 1524 4961 1624 4971
rect 1714 4961 1954 4971
rect 2544 4961 2784 4971
rect 3274 4961 4104 4971
rect 1504 4941 1624 4961
rect 1724 4951 1954 4961
rect 2584 4951 2784 4961
rect 3324 4951 4084 4961
rect 4374 4951 4394 4961
rect 1724 4941 1944 4951
rect 2594 4941 2794 4951
rect 3344 4941 4094 4951
rect 1524 4931 1544 4941
rect 1554 4931 1624 4941
rect 1734 4931 1944 4941
rect 2644 4931 2814 4941
rect 3364 4931 4114 4941
rect 4384 4931 4394 4951
rect 1734 4921 1934 4931
rect 2664 4921 2824 4931
rect 3384 4921 4114 4931
rect 1744 4911 1934 4921
rect 2674 4911 2824 4921
rect 2854 4911 2864 4921
rect 3404 4911 4114 4921
rect 1754 4851 1934 4911
rect 2704 4901 2834 4911
rect 2854 4901 2874 4911
rect 3564 4901 4114 4911
rect 2384 4891 2534 4901
rect 2744 4891 2764 4901
rect 2784 4891 2834 4901
rect 3534 4891 3544 4901
rect 3554 4891 3884 4901
rect 3894 4891 4124 4901
rect 2364 4881 2574 4891
rect 2794 4881 2824 4891
rect 3514 4881 3824 4891
rect 3844 4881 3854 4891
rect 3974 4881 4124 4891
rect 2334 4871 2634 4881
rect 3524 4871 3774 4881
rect 4014 4871 4124 4881
rect 2304 4861 2714 4871
rect 3524 4861 3744 4871
rect 4034 4861 4114 4871
rect 2294 4851 2744 4861
rect 3594 4851 3644 4861
rect 3664 4851 3694 4861
rect 1754 4801 1924 4851
rect 2284 4841 2764 4851
rect 3594 4841 3624 4851
rect 2274 4831 2794 4841
rect 2274 4821 2804 4831
rect 2284 4811 2814 4821
rect 2294 4801 2834 4811
rect 3634 4801 3684 4811
rect 1764 4791 1914 4801
rect 1774 4781 1914 4791
rect 1784 4751 1914 4781
rect 2294 4791 2854 4801
rect 3584 4791 3864 4801
rect 2294 4771 2864 4791
rect 3574 4781 3944 4791
rect 3564 4771 3964 4781
rect 2304 4761 2874 4771
rect 3544 4761 3984 4771
rect 2324 4751 2434 4761
rect 2474 4751 2874 4761
rect 3524 4751 3994 4761
rect 1784 4641 1904 4751
rect 2364 4741 2444 4751
rect 2474 4741 2734 4751
rect 2754 4741 2884 4751
rect 3514 4741 4004 4751
rect 2364 4731 2464 4741
rect 2394 4721 2464 4731
rect 2474 4721 2724 4741
rect 2764 4731 2894 4741
rect 3494 4731 4014 4741
rect 2764 4721 2904 4731
rect 3484 4721 4024 4731
rect 2414 4711 2704 4721
rect 2774 4711 2914 4721
rect 3474 4711 4034 4721
rect 2414 4701 2694 4711
rect 2424 4691 2694 4701
rect 2784 4691 2914 4711
rect 3464 4701 4044 4711
rect 3454 4691 3864 4701
rect 3884 4691 4044 4701
rect 2434 4681 2674 4691
rect 2764 4681 2904 4691
rect 3444 4681 3574 4691
rect 3614 4681 3864 4691
rect 3904 4681 4034 4691
rect 2494 4671 2664 4681
rect 2724 4671 2904 4681
rect 3434 4671 3564 4681
rect 3614 4671 3854 4681
rect 3914 4671 4054 4681
rect 2544 4661 2694 4671
rect 2734 4661 2904 4671
rect 2564 4651 2654 4661
rect 2664 4651 2704 4661
rect 2774 4651 2784 4661
rect 2874 4651 2904 4661
rect 3444 4661 3544 4671
rect 3624 4661 3844 4671
rect 2584 4641 2644 4651
rect 2674 4641 2704 4651
rect 3444 4641 3534 4661
rect 3634 4651 3844 4661
rect 3934 4661 4054 4671
rect 3934 4651 4034 4661
rect 3634 4641 3834 4651
rect 3924 4641 4024 4651
rect 1794 4621 1904 4641
rect 2614 4631 2634 4641
rect 3454 4631 3484 4641
rect 3494 4631 3544 4641
rect 3644 4631 3824 4641
rect 3924 4631 3964 4641
rect 3464 4621 3474 4631
rect 3494 4621 3554 4631
rect 3654 4621 3814 4631
rect 3914 4621 3944 4631
rect 1804 4581 1894 4621
rect 3664 4611 3814 4621
rect 3904 4611 3934 4621
rect 3664 4601 3794 4611
rect 1814 4561 1894 4581
rect 3634 4591 3794 4601
rect 3634 4571 3764 4591
rect 3784 4581 3804 4591
rect 3784 4571 3824 4581
rect 3634 4561 3674 4571
rect 3804 4561 3814 4571
rect 1824 4531 1854 4561
rect 1864 4551 1884 4561
rect 1834 4521 1854 4531
rect 1844 4511 1864 4521
rect 1844 4411 1854 4431
rect 1844 4391 1864 4411
rect 1854 4381 1864 4391
rect 1864 4361 1884 4371
rect 1874 4351 1884 4361
rect 1854 4251 1884 4261
rect 1864 4231 1884 4251
rect 1854 4181 1884 4201
rect 2754 4181 2774 4191
rect 1864 4171 1874 4181
rect 2744 4171 2814 4181
rect 2734 4161 2814 4171
rect 2724 4151 2824 4161
rect 3464 4151 3504 4161
rect 2674 4141 2824 4151
rect 2654 4121 2824 4141
rect 3454 4141 3514 4151
rect 3454 4131 3524 4141
rect 2634 4111 2824 4121
rect 2614 4101 2824 4111
rect 2594 4091 2824 4101
rect 2554 4071 2824 4091
rect 3444 4121 3534 4131
rect 3444 4111 3574 4121
rect 3444 4091 3584 4111
rect 3444 4081 3614 4091
rect 3444 4071 3624 4081
rect 1824 4061 1894 4071
rect 2494 4061 2824 4071
rect 1824 4051 1904 4061
rect 2414 4051 2424 4061
rect 1824 4031 1914 4051
rect 2414 4041 2434 4051
rect 2404 4031 2444 4041
rect 2484 4031 2824 4061
rect 3454 4061 3634 4071
rect 1824 4021 1924 4031
rect 2394 4021 2464 4031
rect 2494 4021 2834 4031
rect 1754 4011 1764 4021
rect 1734 3981 1834 3991
rect 1844 3981 1924 4021
rect 2294 4011 2314 4021
rect 2374 4011 2834 4021
rect 2264 4001 2344 4011
rect 2364 4001 2834 4011
rect 2264 3991 2834 4001
rect 2244 3990 2834 3991
rect 3454 4021 3684 4061
rect 4224 4051 4234 4061
rect 4194 4031 4234 4041
rect 4184 4021 4234 4031
rect 3454 4011 3744 4021
rect 4174 4011 4234 4021
rect 4244 4011 4264 4021
rect 3454 4001 3754 4011
rect 4204 4001 4234 4011
rect 3454 3991 3764 4001
rect 4214 3991 4224 4001
rect 2244 3981 2844 3990
rect 3454 3981 3804 3991
rect 1724 3971 1934 3981
rect 2234 3971 2274 3981
rect 2284 3971 2764 3981
rect 2794 3971 2824 3981
rect 2834 3971 2864 3981
rect 3444 3971 3824 3981
rect 4214 3971 4224 3981
rect 1614 3961 1634 3971
rect 1664 3961 1934 3971
rect 1614 3951 1934 3961
rect 2224 3961 2764 3971
rect 2804 3961 2814 3971
rect 2834 3961 2904 3971
rect 3444 3961 3854 3971
rect 3864 3961 3894 3971
rect 4204 3961 4284 3971
rect 2224 3951 2744 3961
rect 1614 3941 1684 3951
rect 1704 3941 1944 3951
rect 1734 3931 1744 3941
rect 1834 3931 1944 3941
rect 2224 3941 2724 3951
rect 2824 3941 2914 3961
rect 3494 3951 3894 3961
rect 3924 3951 3934 3961
rect 4164 3951 4294 3961
rect 3504 3941 3964 3951
rect 2224 3931 2704 3941
rect 2864 3931 2944 3941
rect 3514 3931 3974 3941
rect 4154 3931 4304 3951
rect 1824 3921 1944 3931
rect 1614 3911 1944 3921
rect 2214 3921 2694 3931
rect 2884 3921 2954 3931
rect 3514 3921 3984 3931
rect 2214 3911 2684 3921
rect 2894 3911 3004 3921
rect 3304 3911 3324 3921
rect 3524 3911 4004 3921
rect 1594 3901 1954 3911
rect 1564 3891 1954 3901
rect 2214 3891 2674 3911
rect 2894 3901 3014 3911
rect 2904 3891 2914 3901
rect 1184 3881 1234 3891
rect 1284 3881 1294 3891
rect 1324 3881 1354 3891
rect 1364 3881 1444 3891
rect 1484 3881 1494 3891
rect 1554 3881 1954 3891
rect 2224 3881 2664 3891
rect 2924 3881 3024 3901
rect 3204 3891 3264 3901
rect 3114 3881 3274 3891
rect 3284 3881 3334 3911
rect 3534 3901 4004 3911
rect 4144 3901 4294 3931
rect 3554 3891 4014 3901
rect 4144 3891 4314 3901
rect 3554 3881 4024 3891
rect 4134 3881 4314 3891
rect 1134 3871 1154 3881
rect 1174 3871 1254 3881
rect 1264 3871 1304 3881
rect 1314 3871 1454 3881
rect 1484 3871 1954 3881
rect 2244 3871 2654 3881
rect 2924 3871 3044 3881
rect 3104 3871 3224 3881
rect 3234 3871 3324 3881
rect 3534 3871 4004 3881
rect 4134 3871 4324 3881
rect 1134 3861 1824 3871
rect 1854 3861 1964 3871
rect 1134 3851 1814 3861
rect 1874 3851 1964 3861
rect 2214 3861 2644 3871
rect 2934 3861 3064 3871
rect 3074 3861 3224 3871
rect 3244 3861 3314 3871
rect 3534 3861 4024 3871
rect 2214 3851 2634 3861
rect 2944 3851 3224 3861
rect 3234 3851 3304 3861
rect 1134 3841 1804 3851
rect 1884 3841 1974 3851
rect 2214 3841 2254 3851
rect 2264 3841 2644 3851
rect 2924 3841 2934 3851
rect 2954 3841 3304 3851
rect 1134 3831 1774 3841
rect 1134 3821 1764 3831
rect 1884 3821 1984 3841
rect 2294 3831 2644 3841
rect 2944 3831 3304 3841
rect 3564 3841 4024 3861
rect 4124 3861 4324 3871
rect 4124 3851 4334 3861
rect 4124 3841 4344 3851
rect 3564 3831 4004 3841
rect 4134 3831 4364 3841
rect 1134 3811 1744 3821
rect 1134 3801 1734 3811
rect 1874 3801 1984 3821
rect 2284 3821 2654 3831
rect 2944 3821 3294 3831
rect 3554 3821 3984 3831
rect 4134 3821 4444 3831
rect 2284 3811 2684 3821
rect 2964 3811 2974 3821
rect 2984 3811 3284 3821
rect 3544 3811 3974 3821
rect 4134 3811 4464 3821
rect 2284 3801 2694 3811
rect 2994 3801 3274 3811
rect 3534 3801 3974 3811
rect 4124 3801 4464 3811
rect 1134 3791 1724 3801
rect 1884 3791 1994 3801
rect 2274 3791 2744 3801
rect 3004 3791 3264 3801
rect 3514 3791 3974 3801
rect 4114 3791 4474 3801
rect 1134 3771 1714 3791
rect 1874 3771 2004 3791
rect 2174 3771 2194 3791
rect 2264 3781 2754 3791
rect 3024 3781 3244 3791
rect 3494 3781 3954 3791
rect 2244 3771 2294 3781
rect 2304 3771 2764 3781
rect 3044 3771 3214 3781
rect 3474 3771 3964 3781
rect 1134 3751 1694 3771
rect 1874 3751 2014 3771
rect 2164 3751 2184 3771
rect 2244 3761 2254 3771
rect 2284 3761 2324 3771
rect 2334 3761 2364 3771
rect 2384 3761 2834 3771
rect 3064 3761 3074 3771
rect 3114 3761 3154 3771
rect 3194 3761 3204 3771
rect 3444 3761 3964 3771
rect 4104 3771 4484 3791
rect 4104 3761 4474 3771
rect 2294 3751 2324 3761
rect 2394 3751 2844 3761
rect 2884 3751 2904 3761
rect 3134 3751 3144 3761
rect 3434 3751 3974 3761
rect 1134 3731 1684 3751
rect 1874 3741 2024 3751
rect 2394 3741 2914 3751
rect 2974 3741 2994 3751
rect 3014 3741 3034 3751
rect 3384 3741 3974 3751
rect 4094 3741 4494 3761
rect 1864 3731 1894 3741
rect 1924 3731 2024 3741
rect 2164 3731 2174 3741
rect 2394 3731 2694 3741
rect 1134 3711 1674 3731
rect 1874 3721 1894 3731
rect 1934 3721 2034 3731
rect 1874 3711 1904 3721
rect 1944 3711 2024 3721
rect 2154 3711 2184 3731
rect 2404 3721 2694 3731
rect 2704 3731 3054 3741
rect 3334 3731 3674 3741
rect 3694 3731 3794 3741
rect 3834 3731 3844 3741
rect 3854 3731 3994 3741
rect 2704 3721 2754 3731
rect 2784 3721 3094 3731
rect 3164 3721 3654 3731
rect 3694 3721 3784 3731
rect 3864 3721 3944 3731
rect 3954 3721 3994 3731
rect 4094 3731 4544 3741
rect 4094 3721 4694 3731
rect 2404 3711 2744 3721
rect 2804 3711 3624 3721
rect 1134 3701 1664 3711
rect 1874 3701 1894 3711
rect 1944 3701 2034 3711
rect 2414 3701 2544 3711
rect 2554 3701 2734 3711
rect 2814 3701 3414 3711
rect 3454 3701 3614 3711
rect 3704 3701 3784 3721
rect 3854 3714 3994 3721
rect 3852 3711 3994 3714
rect 4084 3711 4714 3721
rect 3852 3701 3984 3711
rect 4074 3701 4724 3711
rect 1134 3691 1654 3701
rect 1834 3691 1844 3701
rect 1854 3691 1894 3701
rect 1924 3691 2044 3701
rect 2414 3691 2534 3701
rect 2564 3691 2734 3701
rect 2824 3691 3404 3701
rect 3454 3691 3604 3701
rect 3704 3691 3774 3701
rect 3852 3699 3974 3701
rect 3864 3691 3974 3699
rect 4064 3691 4724 3701
rect 1134 3681 1614 3691
rect 1824 3681 1884 3691
rect 1924 3681 2054 3691
rect 2194 3681 2204 3691
rect 1134 3671 1604 3681
rect 1824 3671 1864 3681
rect 1914 3671 2054 3681
rect 2184 3671 2204 3681
rect 2424 3671 2514 3691
rect 2584 3671 2734 3691
rect 2834 3681 3394 3691
rect 3454 3681 3594 3691
rect 3704 3681 3754 3691
rect 3864 3681 3944 3691
rect 4054 3681 4714 3691
rect 2834 3671 3384 3681
rect 3454 3671 3584 3681
rect 3714 3671 3754 3681
rect 3874 3671 3954 3681
rect 4054 3671 4704 3681
rect 1134 3661 1544 3671
rect 1804 3661 1854 3671
rect 1134 3641 1534 3661
rect 1824 3651 1854 3661
rect 1894 3661 2064 3671
rect 1894 3651 2074 3661
rect 2414 3651 2514 3671
rect 2604 3661 2734 3671
rect 2904 3661 3374 3671
rect 3454 3661 3574 3671
rect 3714 3661 3744 3671
rect 3874 3661 3974 3671
rect 1914 3641 2084 3651
rect 1134 3631 1514 3641
rect 1904 3631 2084 3641
rect 2424 3641 2514 3651
rect 2614 3641 2734 3661
rect 2914 3651 2984 3661
rect 3014 3651 3314 3661
rect 3334 3651 3364 3661
rect 3454 3651 3564 3661
rect 3714 3651 3734 3661
rect 3904 3651 3934 3661
rect 3954 3651 3974 3661
rect 1134 3621 1504 3631
rect 1884 3621 2094 3631
rect 1134 3611 1494 3621
rect 1134 3601 1484 3611
rect 1134 3591 1474 3601
rect 1134 3571 1464 3591
rect 1874 3581 2104 3621
rect 2424 3611 2524 3641
rect 2634 3631 2734 3641
rect 2924 3641 2964 3651
rect 3034 3641 3294 3651
rect 3344 3641 3364 3651
rect 3464 3641 3554 3651
rect 3844 3641 3864 3651
rect 3914 3641 3934 3651
rect 3964 3641 3974 3651
rect 4044 3641 4304 3671
rect 2924 3631 2954 3641
rect 3064 3631 3164 3641
rect 3244 3631 3284 3641
rect 3454 3631 3544 3641
rect 3924 3631 3934 3641
rect 4044 3631 4194 3641
rect 4204 3631 4304 3641
rect 2664 3621 2744 3631
rect 2834 3621 2844 3631
rect 2934 3621 2944 3631
rect 3074 3621 3144 3631
rect 3264 3621 3274 3631
rect 3454 3621 3534 3631
rect 3924 3621 3944 3631
rect 4044 3621 4184 3631
rect 4214 3621 4294 3631
rect 2434 3601 2524 3611
rect 2704 3611 2744 3621
rect 2824 3611 2854 3621
rect 2704 3601 2754 3611
rect 2814 3601 2864 3611
rect 2444 3581 2524 3601
rect 2714 3591 2734 3601
rect 2744 3591 2864 3601
rect 3094 3601 3124 3621
rect 3344 3611 3354 3621
rect 3444 3611 3494 3621
rect 3874 3611 3884 3621
rect 3924 3611 3954 3621
rect 4064 3611 4174 3621
rect 4234 3611 4274 3621
rect 3094 3591 3114 3601
rect 3334 3591 3374 3611
rect 3444 3601 3484 3611
rect 3704 3601 3714 3611
rect 3874 3601 3954 3611
rect 4094 3601 4144 3611
rect 3444 3591 3464 3601
rect 3884 3591 3944 3601
rect 2754 3581 2874 3591
rect 3324 3581 3394 3591
rect 3884 3581 3904 3591
rect 1134 3551 1444 3571
rect 1134 3541 1424 3551
rect 1864 3541 2104 3581
rect 2434 3571 2534 3581
rect 2754 3571 2884 3581
rect 3314 3571 3404 3581
rect 3874 3571 3904 3581
rect 2444 3551 2534 3571
rect 2764 3561 2894 3571
rect 2924 3561 2944 3571
rect 3294 3561 3394 3571
rect 3854 3561 3904 3571
rect 3924 3561 3934 3571
rect 2794 3551 2954 3561
rect 3254 3551 3394 3561
rect 3844 3551 3934 3561
rect 2444 3541 2544 3551
rect 2804 3541 2954 3551
rect 1134 3531 1414 3541
rect 1134 3521 1384 3531
rect 1134 3511 1364 3521
rect 1844 3511 2104 3541
rect 2434 3531 2454 3541
rect 2464 3531 2544 3541
rect 2844 3531 2954 3541
rect 3244 3541 3374 3551
rect 3834 3541 3924 3551
rect 3244 3531 3364 3541
rect 3744 3531 3764 3541
rect 2474 3521 2544 3531
rect 2854 3521 2984 3531
rect 3244 3521 3354 3531
rect 2484 3511 2494 3521
rect 2534 3511 2544 3521
rect 2864 3511 3014 3521
rect 3234 3511 3314 3521
rect 3734 3511 3764 3531
rect 3834 3531 3854 3541
rect 3834 3521 3864 3531
rect 3784 3511 3794 3521
rect 3804 3511 3864 3521
rect 3874 3521 3914 3541
rect 3874 3511 3904 3521
rect 1134 3501 1354 3511
rect 1834 3501 2104 3511
rect 1134 3491 1344 3501
rect 1134 3471 1334 3491
rect 1824 3481 2094 3501
rect 2474 3491 2494 3511
rect 2884 3501 3064 3511
rect 3084 3501 3114 3511
rect 3154 3501 3294 3511
rect 2924 3491 3254 3501
rect 2954 3481 3224 3491
rect 3774 3481 3864 3511
rect 1814 3471 2094 3481
rect 3014 3471 3184 3481
rect 3744 3471 3864 3481
rect 1134 3461 1304 3471
rect 1134 3451 1294 3461
rect 1804 3451 2094 3471
rect 3084 3461 3104 3471
rect 3734 3461 3864 3471
rect 1134 3441 1284 3451
rect 1804 3441 2084 3451
rect 2454 3441 2464 3461
rect 3714 3451 3854 3461
rect 3714 3441 3844 3451
rect 1134 3431 1274 3441
rect 1134 3421 1264 3431
rect 1134 3411 1244 3421
rect 1804 3411 2074 3441
rect 2854 3421 2934 3431
rect 3364 3421 3374 3441
rect 3724 3431 3844 3441
rect 3724 3421 3824 3431
rect 3834 3421 3844 3431
rect 2834 3411 2934 3421
rect 3714 3411 3824 3421
rect 1134 3401 1234 3411
rect 1804 3401 2064 3411
rect 2834 3401 2944 3411
rect 3244 3401 3254 3411
rect 3704 3401 3824 3411
rect 3834 3401 3854 3411
rect 1134 3391 1224 3401
rect 1804 3391 2054 3401
rect 1134 3381 1214 3391
rect 1134 3371 1194 3381
rect 1794 3371 2054 3391
rect 2364 3381 2374 3401
rect 2850 3399 2954 3401
rect 2864 3391 2954 3399
rect 3234 3391 3254 3401
rect 3274 3391 3294 3401
rect 3704 3391 3854 3401
rect 3884 3391 3904 3401
rect 2864 3381 2964 3391
rect 3034 3381 3064 3391
rect 3124 3381 3134 3391
rect 3224 3390 3254 3391
rect 3264 3390 3294 3391
rect 3224 3381 3294 3390
rect 2884 3371 2974 3381
rect 3024 3371 3064 3381
rect 3074 3371 3094 3381
rect 3114 3371 3164 3381
rect 3214 3371 3234 3381
rect 3254 3371 3294 3381
rect 3694 3381 3854 3391
rect 3874 3381 3904 3391
rect 3694 3371 3864 3381
rect 1134 3351 1184 3371
rect 1784 3361 2054 3371
rect 2894 3361 2904 3371
rect 2914 3361 2984 3371
rect 2994 3361 3104 3371
rect 3114 3361 3284 3371
rect 3304 3361 3324 3371
rect 3704 3361 3864 3371
rect 1784 3351 2044 3361
rect 1134 3341 1174 3351
rect 1144 3331 1154 3341
rect 1774 3311 2034 3351
rect 2344 3331 2364 3341
rect 2334 3321 2364 3331
rect 2924 3331 3324 3361
rect 3384 3341 3404 3361
rect 3674 3341 3894 3361
rect 3374 3331 3394 3341
rect 3664 3331 3894 3341
rect 2924 3321 2954 3331
rect 2344 3311 2374 3321
rect 2824 3311 2844 3321
rect 2914 3311 2954 3321
rect 2964 3321 3324 3331
rect 3344 3321 3384 3331
rect 3664 3321 3904 3331
rect 2964 3311 3374 3321
rect 1774 3301 2024 3311
rect 2354 3301 2364 3311
rect 2424 3301 2444 3311
rect 1764 3291 2024 3301
rect 2414 3291 2444 3301
rect 2814 3301 2844 3311
rect 2864 3301 2874 3311
rect 2904 3301 3374 3311
rect 3654 3301 3914 3321
rect 2814 3291 2834 3301
rect 2864 3291 3364 3301
rect 3634 3291 3914 3301
rect 1754 3261 2014 3291
rect 2344 3271 2444 3291
rect 2764 3281 2784 3291
rect 2824 3281 2834 3291
rect 2884 3281 3354 3291
rect 3624 3281 3924 3291
rect 2884 3271 3324 3281
rect 3624 3271 3934 3281
rect 2344 3261 2404 3271
rect 2424 3261 2444 3271
rect 2874 3261 3324 3271
rect 3614 3261 3944 3271
rect 1754 3241 2004 3261
rect 2344 3251 2434 3261
rect 2454 3251 2464 3261
rect 2884 3251 3314 3261
rect 3604 3251 3924 3261
rect 3934 3251 3944 3261
rect 1744 3231 2004 3241
rect 2384 3231 2424 3251
rect 2454 3241 2474 3251
rect 2894 3241 3254 3251
rect 3264 3241 3294 3251
rect 2454 3231 2504 3241
rect 2914 3231 2934 3241
rect 2984 3231 3254 3241
rect 1734 3211 2004 3231
rect 2394 3221 2424 3231
rect 2464 3221 2514 3231
rect 3004 3221 3084 3231
rect 3124 3221 3134 3231
rect 3244 3221 3254 3231
rect 3584 3221 3904 3251
rect 2394 3211 2454 3221
rect 2474 3211 2514 3221
rect 3054 3211 3074 3221
rect 3574 3211 3914 3221
rect 1744 3191 1994 3211
rect 2404 3201 2454 3211
rect 2484 3201 2494 3211
rect 1734 3181 1994 3191
rect 2364 3183 2394 3192
rect 2414 3191 2474 3201
rect 3564 3191 3924 3211
rect 2364 3181 2385 3183
rect 2414 3181 2554 3191
rect 3564 3181 3914 3191
rect 1734 3171 1984 3181
rect 2374 3171 2385 3181
rect 2404 3171 2554 3181
rect 3554 3171 3924 3181
rect 1734 3161 1974 3171
rect 2394 3161 2564 3171
rect 3544 3161 3934 3171
rect 1724 3141 1974 3161
rect 1714 3131 1974 3141
rect 2404 3151 2564 3161
rect 3534 3151 3934 3161
rect 2404 3141 2574 3151
rect 2404 3131 2594 3141
rect 3534 3131 3944 3151
rect 1724 3121 1964 3131
rect 2424 3121 2604 3131
rect 3534 3121 3934 3131
rect 1724 3111 1954 3121
rect 1714 3101 1954 3111
rect 1704 3071 1954 3101
rect 2434 3111 2604 3121
rect 3514 3111 3934 3121
rect 2434 3091 2614 3111
rect 3504 3101 3924 3111
rect 2424 3081 2634 3091
rect 3504 3081 3934 3101
rect 2424 3071 2644 3081
rect 3494 3071 3934 3081
rect 1714 3061 1954 3071
rect 2454 3061 2654 3071
rect 1714 3041 1944 3061
rect 2434 3045 2444 3051
rect 2464 3045 2654 3061
rect 3484 3061 3964 3071
rect 3484 3051 3954 3061
rect 2434 3041 2654 3045
rect 3454 3041 3464 3051
rect 3474 3041 3954 3051
rect 1714 3031 1954 3041
rect 2434 3031 2674 3041
rect 3444 3031 3954 3041
rect 1704 3001 1934 3031
rect 2442 3030 2694 3031
rect 2454 3021 2694 3030
rect 3434 3021 3954 3031
rect 2444 3011 2704 3021
rect 3424 3011 3964 3021
rect 2454 3001 2464 3011
rect 2484 3001 2714 3011
rect 3394 3001 3974 3011
rect 1684 2961 1934 3001
rect 2484 2991 2724 3001
rect 2734 2991 2744 3001
rect 3374 2991 3974 3001
rect 2494 2981 2764 2991
rect 3364 2981 3974 2991
rect 2534 2971 2774 2981
rect 3334 2971 3984 2981
rect 2464 2961 2514 2971
rect 2534 2961 2804 2971
rect 3294 2961 3974 2971
rect 1684 2951 1924 2961
rect 2454 2951 2824 2961
rect 3284 2951 3974 2961
rect 1684 2941 1934 2951
rect 2474 2941 2844 2951
rect 2874 2941 2894 2951
rect 2924 2941 2944 2951
rect 2954 2941 2984 2951
rect 3004 2941 3074 2951
rect 3104 2941 3174 2951
rect 3204 2941 3974 2951
rect 1674 2871 1934 2941
rect 2484 2921 2894 2941
rect 2914 2931 3074 2941
rect 3094 2931 3964 2941
rect 2904 2921 3074 2931
rect 3084 2921 3964 2931
rect 2504 2911 3964 2921
rect 2454 2891 2464 2911
rect 2514 2901 3964 2911
rect 2514 2891 3974 2901
rect 2474 2881 2554 2891
rect 2564 2881 3974 2891
rect 2484 2871 2534 2881
rect 2574 2871 3974 2881
rect 1664 2861 1934 2871
rect 2494 2861 2524 2871
rect 2564 2861 3984 2871
rect 1664 2841 1944 2861
rect 2534 2851 3984 2861
rect 2394 2841 2434 2851
rect 2544 2841 3984 2851
rect 1654 2821 1924 2841
rect 2404 2831 2444 2841
rect 2354 2821 2364 2831
rect 2414 2821 2454 2831
rect 2594 2821 3984 2841
rect 1654 2811 1934 2821
rect 2344 2811 2374 2821
rect 2424 2811 2454 2821
rect 2534 2811 3984 2821
rect 1654 2771 1944 2811
rect 2424 2801 2514 2811
rect 2524 2801 3984 2811
rect 2424 2791 3984 2801
rect 2304 2781 2324 2791
rect 2424 2781 2504 2791
rect 2524 2781 3984 2791
rect 2294 2771 2334 2781
rect 2384 2771 2414 2781
rect 2434 2771 2484 2781
rect 2534 2771 3984 2781
rect 1654 2761 1954 2771
rect 2324 2761 2344 2771
rect 2544 2761 3984 2771
rect 4004 2761 4014 2781
rect 1654 2741 1944 2761
rect 2324 2741 2354 2761
rect 2454 2751 2474 2761
rect 2544 2751 4014 2761
rect 2424 2741 2484 2751
rect 1654 2731 1934 2741
rect 1644 2701 1944 2731
rect 2264 2721 2284 2741
rect 2324 2731 2344 2741
rect 2434 2731 2494 2741
rect 2534 2731 2634 2751
rect 2664 2741 4014 2751
rect 2654 2731 4014 2741
rect 2314 2721 2344 2731
rect 2394 2721 2414 2731
rect 2434 2721 2514 2731
rect 2314 2711 2334 2721
rect 2404 2711 2424 2721
rect 2474 2711 2504 2721
rect 2544 2711 4024 2731
rect 2304 2701 2354 2711
rect 2414 2701 2494 2711
rect 2534 2701 4034 2711
rect 1644 2681 1954 2701
rect 2304 2691 2364 2701
rect 2414 2691 4024 2701
rect 2264 2681 2294 2691
rect 2314 2681 2354 2691
rect 2414 2682 2544 2691
rect 1634 2671 1954 2681
rect 2314 2671 2344 2681
rect 2412 2671 2544 2682
rect 2554 2681 4034 2691
rect 2564 2671 4044 2681
rect 1634 2661 1944 2671
rect 2314 2661 2374 2671
rect 2412 2670 2436 2671
rect 2414 2661 2424 2670
rect 2464 2661 4054 2671
rect 1624 2651 1934 2661
rect 2234 2651 2254 2661
rect 2304 2651 2374 2661
rect 2404 2651 2424 2661
rect 2454 2651 4054 2661
rect 1624 2641 1954 2651
rect 1634 2621 1954 2641
rect 2224 2641 2264 2651
rect 2314 2641 2484 2651
rect 2504 2641 4054 2651
rect 2224 2631 2254 2641
rect 2324 2631 4054 2641
rect 2224 2621 2244 2631
rect 1634 2611 1934 2621
rect 2294 2611 2314 2631
rect 2334 2621 4064 2631
rect 2364 2611 4064 2621
rect 1624 2601 1934 2611
rect 2244 2601 2264 2611
rect 1624 2581 1884 2601
rect 2234 2591 2264 2601
rect 2304 2591 4074 2611
rect 1944 2581 1964 2591
rect 2244 2581 2264 2591
rect 2284 2581 2404 2591
rect 2414 2581 4084 2591
rect 1624 2571 1894 2581
rect 1944 2571 1974 2581
rect 2284 2571 4094 2581
rect 1624 2551 1914 2571
rect 2284 2561 2314 2571
rect 2334 2561 4104 2571
rect 2334 2551 4114 2561
rect 1624 2541 1874 2551
rect 2264 2541 2284 2551
rect 2334 2541 4074 2551
rect 4094 2541 4114 2551
rect 1624 2521 1884 2541
rect 2194 2531 2234 2541
rect 2204 2521 2234 2531
rect 2264 2521 2294 2541
rect 2344 2531 4064 2541
rect 1624 2511 1854 2521
rect 2314 2511 2324 2521
rect 2354 2511 4044 2531
rect 1624 2501 1864 2511
rect 1624 2491 1854 2501
rect 2304 2491 4044 2511
rect 4414 2511 4424 2521
rect 4414 2491 4434 2511
rect 1624 2481 1834 2491
rect 2324 2481 4044 2491
rect 1614 2471 1834 2481
rect 2124 2471 2144 2481
rect 1614 2461 1814 2471
rect 2224 2461 2254 2471
rect 2334 2461 2354 2481
rect 2364 2461 4054 2481
rect 1624 2451 1814 2461
rect 2214 2451 2264 2461
rect 1624 2431 1824 2451
rect 2234 2441 2264 2451
rect 2294 2441 2324 2461
rect 2334 2441 4054 2461
rect 2124 2431 2144 2441
rect 2244 2431 2254 2441
rect 1624 2421 1814 2431
rect 1624 2401 1804 2421
rect 2244 2411 2254 2421
rect 2344 2411 2374 2441
rect 2394 2431 4064 2441
rect 4334 2431 4344 2441
rect 4424 2431 4444 2441
rect 2384 2411 4074 2431
rect 4334 2421 4364 2431
rect 4414 2421 4494 2431
rect 4324 2411 4374 2421
rect 4404 2411 4494 2421
rect 2234 2401 2264 2411
rect 2294 2401 2314 2411
rect 2344 2401 4084 2411
rect 4304 2401 4484 2411
rect 1624 2381 1784 2401
rect 2294 2391 2324 2401
rect 2354 2391 2374 2401
rect 2384 2391 2404 2401
rect 2304 2381 2324 2391
rect 2424 2381 4084 2401
rect 4294 2391 4394 2401
rect 4414 2391 4444 2401
rect 4454 2391 4484 2401
rect 4294 2381 4384 2391
rect 4464 2381 4484 2391
rect 1624 2371 1764 2381
rect 2384 2371 2394 2381
rect 2434 2371 4094 2381
rect 4304 2371 4414 2381
rect 1624 2361 1754 2371
rect 2314 2361 2334 2371
rect 1624 2341 1744 2361
rect 2324 2351 2334 2361
rect 2354 2361 4094 2371
rect 4314 2361 4434 2371
rect 2354 2351 2424 2361
rect 1764 2341 1774 2351
rect 2374 2341 2424 2351
rect 2454 2351 4104 2361
rect 4324 2351 4454 2361
rect 4464 2351 4494 2361
rect 2454 2341 2514 2351
rect 2524 2341 4104 2351
rect 4334 2341 4494 2351
rect 1624 2331 1774 2341
rect 2334 2331 2354 2341
rect 2464 2331 2504 2341
rect 2554 2331 4104 2341
rect 4364 2331 4524 2341
rect 1624 2311 1744 2331
rect 2374 2321 2394 2331
rect 1614 2301 1744 2311
rect 2364 2301 2404 2321
rect 2454 2311 2514 2331
rect 2534 2321 4114 2331
rect 4394 2321 4524 2331
rect 2534 2311 2564 2321
rect 2594 2311 2634 2321
rect 2454 2301 2504 2311
rect 2544 2301 2564 2311
rect 2604 2301 2634 2311
rect 2644 2311 4114 2321
rect 4414 2311 4554 2321
rect 2644 2301 4124 2311
rect 4424 2301 4584 2311
rect 1614 2281 1734 2301
rect 2374 2291 2394 2301
rect 2384 2281 2394 2291
rect 2464 2281 2494 2301
rect 2584 2291 3344 2301
rect 3354 2291 4124 2301
rect 4454 2291 4584 2301
rect 2584 2281 2654 2291
rect 2674 2281 3344 2291
rect 3364 2281 4124 2291
rect 4464 2281 4594 2291
rect 1134 2271 1154 2281
rect 1614 2271 1724 2281
rect 2454 2271 2494 2281
rect 2595 2280 2646 2281
rect 1134 2241 1174 2271
rect 1614 2251 1734 2271
rect 2464 2261 2484 2271
rect 2604 2261 2634 2280
rect 2674 2271 4124 2281
rect 4504 2271 4594 2281
rect 2654 2261 3374 2271
rect 3384 2261 4134 2271
rect 4514 2261 4604 2271
rect 4634 2261 4654 2271
rect 2644 2251 2684 2261
rect 2744 2251 2784 2261
rect 2794 2251 3204 2261
rect 1144 2231 1174 2241
rect 1624 2231 1724 2251
rect 2644 2241 2674 2251
rect 2754 2241 2784 2251
rect 2814 2241 2834 2251
rect 2854 2241 2934 2251
rect 2954 2241 3134 2251
rect 3154 2241 3204 2251
rect 3234 2251 4134 2261
rect 4554 2251 4664 2261
rect 3234 2241 3274 2251
rect 3284 2250 4144 2251
rect 2514 2231 2534 2241
rect 2564 2231 2584 2241
rect 2704 2231 2734 2241
rect 2864 2231 2914 2241
rect 2964 2231 3273 2241
rect 3284 2231 3304 2250
rect 3314 2241 4144 2250
rect 4564 2241 4664 2251
rect 3344 2231 4154 2241
rect 4574 2231 4664 2241
rect 1614 2211 1714 2231
rect 2504 2221 2534 2231
rect 2554 2221 2584 2231
rect 2604 2221 2614 2231
rect 2654 2221 2714 2231
rect 2884 2221 2904 2231
rect 3004 2221 3054 2231
rect 2564 2211 2574 2221
rect 2654 2211 2694 2221
rect 3014 2211 3054 2221
rect 3094 2221 3156 2231
rect 3204 2229 3314 2231
rect 3204 2221 3254 2229
rect 3094 2211 3164 2221
rect 3214 2211 3244 2221
rect 3264 2211 3314 2229
rect 3364 2221 4154 2231
rect 4594 2221 4654 2231
rect 1604 2181 1714 2211
rect 2534 2201 2544 2211
rect 2534 2191 2554 2201
rect 3024 2191 3054 2211
rect 3144 2201 3164 2211
rect 3364 2201 4164 2221
rect 4624 2211 4654 2221
rect 2534 2181 2574 2191
rect 1614 2161 1724 2181
rect 2974 2171 2984 2191
rect 3034 2181 3054 2191
rect 3084 2191 3104 2201
rect 3354 2191 4174 2201
rect 3084 2181 3094 2191
rect 3344 2171 4174 2191
rect 3154 2161 3194 2171
rect 3344 2161 4184 2171
rect 1624 2141 1734 2161
rect 3114 2151 3124 2161
rect 3364 2151 4184 2161
rect 3364 2141 4194 2151
rect 1634 2131 1724 2141
rect 3324 2131 4194 2141
rect 1624 2121 1724 2131
rect 3314 2121 4204 2131
rect 1614 2111 1734 2121
rect 1624 2071 1734 2111
rect 3324 2091 4204 2121
rect 1744 2071 1764 2081
rect 1624 2021 1764 2071
rect 3324 2051 4224 2091
rect 3314 2041 4234 2051
rect 3314 2031 4244 2041
rect 1624 2001 1774 2021
rect 3304 2001 4244 2031
rect 1634 1981 1774 2001
rect 3284 1981 4244 2001
rect 1624 1961 1774 1981
rect 3274 1971 4254 1981
rect 3274 1961 4264 1971
rect 1634 1931 1784 1961
rect 3284 1941 4264 1961
rect 3294 1931 4274 1941
rect 1624 1911 1784 1931
rect 3274 1921 4274 1931
rect 1624 1901 1774 1911
rect 3254 1901 4274 1921
rect 1624 1891 1764 1901
rect 3244 1891 4284 1901
rect 1614 1871 1764 1891
rect 3234 1881 4284 1891
rect 3234 1871 4294 1881
rect 1604 1841 1764 1871
rect 3244 1861 4294 1871
rect 1594 1821 1764 1841
rect 3234 1851 4294 1861
rect 3234 1831 4304 1851
rect 1584 1811 1764 1821
rect 3224 1821 4304 1831
rect 1574 1801 1754 1811
rect 3224 1801 4314 1821
rect 1514 1791 1534 1801
rect 1504 1761 1544 1791
rect 1414 1741 1444 1761
rect 1494 1751 1534 1761
rect 1484 1741 1524 1751
rect 1474 1731 1514 1741
rect 1464 1721 1514 1731
rect 1464 1711 1504 1721
rect 1454 1701 1494 1711
rect 1444 1691 1484 1701
rect 1364 1681 1394 1691
rect 1354 1661 1394 1681
rect 1434 1681 1474 1691
rect 1434 1671 1464 1681
rect 1434 1661 1444 1671
rect 1354 1651 1404 1661
rect 1574 1651 1734 1801
rect 3224 1791 4324 1801
rect 3214 1761 4324 1791
rect 3204 1741 4334 1761
rect 3174 1731 4344 1741
rect 3164 1711 4344 1731
rect 3154 1691 4344 1711
rect 3154 1671 4354 1691
rect 3144 1661 4364 1671
rect 3124 1651 4364 1661
rect 1354 1641 1384 1651
rect 1334 1621 1384 1641
rect 1324 1611 1384 1621
rect 1574 1611 1714 1651
rect 3114 1641 4374 1651
rect 3104 1631 4374 1641
rect 3094 1611 4374 1631
rect 1314 1591 1334 1611
rect 1354 1601 1384 1611
rect 1354 1591 1374 1601
rect 1324 1581 1364 1591
rect 1264 1571 1294 1581
rect 1324 1571 1354 1581
rect 1254 1561 1294 1571
rect 1564 1561 1714 1611
rect 3084 1591 4384 1611
rect 3074 1581 4394 1591
rect 3054 1561 4394 1581
rect 1244 1551 1324 1561
rect 1244 1541 1314 1551
rect 1244 1531 1304 1541
rect 1564 1531 1704 1561
rect 3054 1541 4404 1561
rect 3034 1531 4404 1541
rect 1254 1521 1284 1531
rect 1564 1521 1714 1531
rect 3024 1521 4414 1531
rect 1254 1511 1274 1521
rect 1174 1501 1184 1511
rect 1214 1501 1224 1511
rect 1164 1491 1194 1501
rect 1154 1481 1194 1491
rect 1564 1491 1724 1521
rect 3014 1511 4414 1521
rect 2994 1501 4414 1511
rect 2974 1491 4424 1501
rect 1564 1471 1734 1491
rect 2974 1481 4434 1491
rect 1554 1431 1734 1471
rect 2994 1461 4434 1481
rect 2974 1441 4444 1461
rect 2944 1431 4444 1441
rect 1554 1421 1744 1431
rect 1554 1401 1754 1421
rect 2934 1411 4454 1431
rect 1554 1341 1764 1401
rect 2934 1391 4464 1411
rect 2904 1381 4464 1391
rect 2874 1371 4464 1381
rect 2874 1361 4474 1371
rect 2884 1341 4474 1361
rect 1554 1331 1804 1341
rect 2874 1331 4484 1341
rect 1554 1311 1794 1331
rect 2874 1321 4494 1331
rect 1554 1301 1804 1311
rect 2864 1301 4494 1321
rect 1554 1291 1814 1301
rect 2854 1291 4494 1301
rect 1554 1261 1824 1291
rect 2844 1281 4504 1291
rect 2834 1271 4504 1281
rect 1554 1251 1814 1261
rect 2824 1251 4514 1271
rect 1554 1241 1824 1251
rect 2814 1241 4524 1251
rect 1554 1221 1834 1241
rect 2754 1221 2774 1231
rect 2794 1221 4524 1241
rect 1564 1212 1874 1221
rect 1564 1201 1893 1212
rect 2744 1211 4534 1221
rect 2734 1201 4534 1211
rect 1564 1200 1904 1201
rect 1564 1191 1864 1200
rect 1884 1191 1904 1200
rect 2714 1191 4534 1201
rect 1554 1181 1904 1191
rect 2704 1181 4524 1191
rect 1554 1171 1884 1181
rect 2694 1171 4514 1181
rect 1564 1141 1884 1171
rect 2684 1161 4514 1171
rect 2664 1151 4504 1161
rect 2654 1141 4504 1151
rect 1564 1131 1914 1141
rect 2654 1131 4494 1141
rect 1564 1121 1934 1131
rect 1564 1091 1954 1121
rect 2644 1111 4494 1131
rect 2634 1101 4484 1111
rect 2614 1091 4494 1101
rect 1564 1081 1944 1091
rect 2594 1081 4494 1091
rect 1564 1071 1964 1081
rect 2584 1071 4494 1081
rect 1564 1041 1984 1071
rect 2574 1061 4504 1071
rect 2544 1051 4504 1061
rect 2034 1041 2044 1051
rect 2534 1041 4514 1051
rect 1554 1031 1994 1041
rect 2534 1031 4524 1041
rect 1554 1021 2004 1031
rect 2524 1021 4524 1031
rect 1554 1011 2024 1021
rect 2484 1011 4524 1021
rect 1554 1001 2054 1011
rect 2474 1001 4524 1011
rect 1554 991 2074 1001
rect 2334 991 2364 1001
rect 2414 991 4524 1001
rect 1554 981 2104 991
rect 1554 971 2134 981
rect 2254 971 2284 981
rect 2314 971 2374 991
rect 2404 981 4534 991
rect 2394 971 4544 981
rect 1554 961 2174 971
rect 2254 961 2294 971
rect 2304 961 4544 971
rect 1554 951 2184 961
rect 2264 951 4544 961
rect 1554 931 4534 951
rect 1554 911 4564 931
rect 1554 901 4574 911
rect 1554 861 4584 901
rect 1554 831 4594 861
rect 1554 821 4604 831
rect 1544 801 4614 821
rect 1544 781 4624 801
rect 1544 741 4634 781
rect 1544 718 4644 741
<< end >>
