magic
tech scmos
timestamp 1259953556
<< nwell >>
rect 4639 152 4683 190
rect 4695 152 4739 190
<< electrodecontact >>
rect 539 125 543 129
rect 545 125 549 129
rect 551 125 555 129
rect 557 125 561 129
rect 563 125 567 129
rect 569 125 573 129
rect 575 125 579 129
rect 539 112 543 116
rect 545 112 549 116
rect 551 112 555 116
rect 557 112 561 116
rect 563 112 567 116
rect 569 112 573 116
rect 575 112 579 116
rect 629 125 633 129
rect 635 125 639 129
rect 641 125 645 129
rect 647 125 651 129
rect 653 125 657 129
rect 659 125 663 129
rect 665 125 669 129
rect 629 112 633 116
rect 635 112 639 116
rect 641 112 645 116
rect 647 112 651 116
rect 653 112 657 116
rect 659 112 663 116
rect 665 112 669 116
rect 540 95 544 99
rect 546 95 550 99
rect 552 95 556 99
rect 558 95 562 99
rect 564 95 568 99
rect 540 89 544 93
rect 546 89 550 93
rect 552 89 556 93
rect 558 89 562 93
rect 564 89 568 93
rect 540 82 544 86
rect 546 82 550 86
rect 552 82 556 86
rect 558 82 562 86
rect 564 82 568 86
rect 540 76 544 80
rect 546 76 550 80
rect 552 76 556 80
rect 558 76 562 80
rect 564 76 568 80
rect 540 70 544 74
rect 546 70 550 74
rect 552 70 556 74
rect 558 70 562 74
rect 564 70 568 74
rect 540 64 544 68
rect 546 64 550 68
rect 552 64 556 68
rect 558 64 562 68
rect 564 64 568 68
rect 640 95 644 99
rect 646 95 650 99
rect 652 95 656 99
rect 658 95 662 99
rect 664 95 668 99
rect 640 89 644 93
rect 646 89 650 93
rect 652 89 656 93
rect 658 89 662 93
rect 664 89 668 93
rect 640 82 644 86
rect 646 82 650 86
rect 652 82 656 86
rect 658 82 662 86
rect 664 82 668 86
rect 640 76 644 80
rect 646 76 650 80
rect 652 76 656 80
rect 658 76 662 80
rect 664 76 668 80
rect 640 70 644 74
rect 646 70 650 74
rect 652 70 656 74
rect 658 70 662 74
rect 664 70 668 74
rect 640 64 644 68
rect 646 64 650 68
rect 652 64 656 68
rect 658 64 662 68
rect 664 64 668 68
rect 573 53 577 57
rect 583 53 587 57
rect 539 38 543 42
rect 545 38 549 42
rect 551 38 555 42
rect 557 38 561 42
rect 563 38 567 42
rect 569 38 573 42
rect 575 38 579 42
rect 539 20 543 24
rect 545 20 549 24
rect 551 20 555 24
rect 557 20 561 24
rect 563 20 567 24
rect 569 20 573 24
rect 575 20 579 24
rect 621 53 625 57
rect 631 53 635 57
rect 629 38 633 42
rect 635 38 639 42
rect 641 38 645 42
rect 647 38 651 42
rect 653 38 657 42
rect 659 38 663 42
rect 665 38 669 42
rect 629 20 633 24
rect 635 20 639 24
rect 641 20 645 24
rect 647 20 651 24
rect 653 20 657 24
rect 659 20 663 24
rect 665 20 669 24
rect 1013 125 1017 129
rect 1019 125 1023 129
rect 1025 125 1029 129
rect 1031 125 1035 129
rect 1037 125 1041 129
rect 1043 125 1047 129
rect 1049 125 1053 129
rect 1013 112 1017 116
rect 1019 112 1023 116
rect 1025 112 1029 116
rect 1031 112 1035 116
rect 1037 112 1041 116
rect 1043 112 1047 116
rect 1049 112 1053 116
rect 1103 125 1107 129
rect 1109 125 1113 129
rect 1115 125 1119 129
rect 1121 125 1125 129
rect 1127 125 1131 129
rect 1133 125 1137 129
rect 1139 125 1143 129
rect 1103 112 1107 116
rect 1109 112 1113 116
rect 1115 112 1119 116
rect 1121 112 1125 116
rect 1127 112 1131 116
rect 1133 112 1137 116
rect 1139 112 1143 116
rect 1014 95 1018 99
rect 1020 95 1024 99
rect 1026 95 1030 99
rect 1032 95 1036 99
rect 1038 95 1042 99
rect 1014 89 1018 93
rect 1020 89 1024 93
rect 1026 89 1030 93
rect 1032 89 1036 93
rect 1038 89 1042 93
rect 1014 82 1018 86
rect 1020 82 1024 86
rect 1026 82 1030 86
rect 1032 82 1036 86
rect 1038 82 1042 86
rect 1014 76 1018 80
rect 1020 76 1024 80
rect 1026 76 1030 80
rect 1032 76 1036 80
rect 1038 76 1042 80
rect 1014 70 1018 74
rect 1020 70 1024 74
rect 1026 70 1030 74
rect 1032 70 1036 74
rect 1038 70 1042 74
rect 1014 64 1018 68
rect 1020 64 1024 68
rect 1026 64 1030 68
rect 1032 64 1036 68
rect 1038 64 1042 68
rect 1114 95 1118 99
rect 1120 95 1124 99
rect 1126 95 1130 99
rect 1132 95 1136 99
rect 1138 95 1142 99
rect 1114 89 1118 93
rect 1120 89 1124 93
rect 1126 89 1130 93
rect 1132 89 1136 93
rect 1138 89 1142 93
rect 1114 82 1118 86
rect 1120 82 1124 86
rect 1126 82 1130 86
rect 1132 82 1136 86
rect 1138 82 1142 86
rect 1114 76 1118 80
rect 1120 76 1124 80
rect 1126 76 1130 80
rect 1132 76 1136 80
rect 1138 76 1142 80
rect 1114 70 1118 74
rect 1120 70 1124 74
rect 1126 70 1130 74
rect 1132 70 1136 74
rect 1138 70 1142 74
rect 1114 64 1118 68
rect 1120 64 1124 68
rect 1126 64 1130 68
rect 1132 64 1136 68
rect 1138 64 1142 68
rect 1047 53 1051 57
rect 1057 53 1061 57
rect 1013 38 1017 42
rect 1019 38 1023 42
rect 1025 38 1029 42
rect 1031 38 1035 42
rect 1037 38 1041 42
rect 1043 38 1047 42
rect 1049 38 1053 42
rect 1013 20 1017 24
rect 1019 20 1023 24
rect 1025 20 1029 24
rect 1031 20 1035 24
rect 1037 20 1041 24
rect 1043 20 1047 24
rect 1049 20 1053 24
rect 1095 53 1099 57
rect 1105 53 1109 57
rect 1103 38 1107 42
rect 1109 38 1113 42
rect 1115 38 1119 42
rect 1121 38 1125 42
rect 1127 38 1131 42
rect 1133 38 1137 42
rect 1139 38 1143 42
rect 1103 20 1107 24
rect 1109 20 1113 24
rect 1115 20 1119 24
rect 1121 20 1125 24
rect 1127 20 1131 24
rect 1133 20 1137 24
rect 1139 20 1143 24
rect 1487 125 1491 129
rect 1493 125 1497 129
rect 1499 125 1503 129
rect 1505 125 1509 129
rect 1511 125 1515 129
rect 1517 125 1521 129
rect 1523 125 1527 129
rect 1487 112 1491 116
rect 1493 112 1497 116
rect 1499 112 1503 116
rect 1505 112 1509 116
rect 1511 112 1515 116
rect 1517 112 1521 116
rect 1523 112 1527 116
rect 1577 125 1581 129
rect 1583 125 1587 129
rect 1589 125 1593 129
rect 1595 125 1599 129
rect 1601 125 1605 129
rect 1607 125 1611 129
rect 1613 125 1617 129
rect 1577 112 1581 116
rect 1583 112 1587 116
rect 1589 112 1593 116
rect 1595 112 1599 116
rect 1601 112 1605 116
rect 1607 112 1611 116
rect 1613 112 1617 116
rect 1488 95 1492 99
rect 1494 95 1498 99
rect 1500 95 1504 99
rect 1506 95 1510 99
rect 1512 95 1516 99
rect 1488 89 1492 93
rect 1494 89 1498 93
rect 1500 89 1504 93
rect 1506 89 1510 93
rect 1512 89 1516 93
rect 1488 82 1492 86
rect 1494 82 1498 86
rect 1500 82 1504 86
rect 1506 82 1510 86
rect 1512 82 1516 86
rect 1488 76 1492 80
rect 1494 76 1498 80
rect 1500 76 1504 80
rect 1506 76 1510 80
rect 1512 76 1516 80
rect 1488 70 1492 74
rect 1494 70 1498 74
rect 1500 70 1504 74
rect 1506 70 1510 74
rect 1512 70 1516 74
rect 1488 64 1492 68
rect 1494 64 1498 68
rect 1500 64 1504 68
rect 1506 64 1510 68
rect 1512 64 1516 68
rect 1588 95 1592 99
rect 1594 95 1598 99
rect 1600 95 1604 99
rect 1606 95 1610 99
rect 1612 95 1616 99
rect 1588 89 1592 93
rect 1594 89 1598 93
rect 1600 89 1604 93
rect 1606 89 1610 93
rect 1612 89 1616 93
rect 1588 82 1592 86
rect 1594 82 1598 86
rect 1600 82 1604 86
rect 1606 82 1610 86
rect 1612 82 1616 86
rect 1588 76 1592 80
rect 1594 76 1598 80
rect 1600 76 1604 80
rect 1606 76 1610 80
rect 1612 76 1616 80
rect 1588 70 1592 74
rect 1594 70 1598 74
rect 1600 70 1604 74
rect 1606 70 1610 74
rect 1612 70 1616 74
rect 1588 64 1592 68
rect 1594 64 1598 68
rect 1600 64 1604 68
rect 1606 64 1610 68
rect 1612 64 1616 68
rect 1521 53 1525 57
rect 1531 53 1535 57
rect 1487 38 1491 42
rect 1493 38 1497 42
rect 1499 38 1503 42
rect 1505 38 1509 42
rect 1511 38 1515 42
rect 1517 38 1521 42
rect 1523 38 1527 42
rect 1487 20 1491 24
rect 1493 20 1497 24
rect 1499 20 1503 24
rect 1505 20 1509 24
rect 1511 20 1515 24
rect 1517 20 1521 24
rect 1523 20 1527 24
rect 1569 53 1573 57
rect 1579 53 1583 57
rect 1577 38 1581 42
rect 1583 38 1587 42
rect 1589 38 1593 42
rect 1595 38 1599 42
rect 1601 38 1605 42
rect 1607 38 1611 42
rect 1613 38 1617 42
rect 1577 20 1581 24
rect 1583 20 1587 24
rect 1589 20 1593 24
rect 1595 20 1599 24
rect 1601 20 1605 24
rect 1607 20 1611 24
rect 1613 20 1617 24
rect 1961 125 1965 129
rect 1967 125 1971 129
rect 1973 125 1977 129
rect 1979 125 1983 129
rect 1985 125 1989 129
rect 1991 125 1995 129
rect 1997 125 2001 129
rect 1961 112 1965 116
rect 1967 112 1971 116
rect 1973 112 1977 116
rect 1979 112 1983 116
rect 1985 112 1989 116
rect 1991 112 1995 116
rect 1997 112 2001 116
rect 2051 125 2055 129
rect 2057 125 2061 129
rect 2063 125 2067 129
rect 2069 125 2073 129
rect 2075 125 2079 129
rect 2081 125 2085 129
rect 2087 125 2091 129
rect 2051 112 2055 116
rect 2057 112 2061 116
rect 2063 112 2067 116
rect 2069 112 2073 116
rect 2075 112 2079 116
rect 2081 112 2085 116
rect 2087 112 2091 116
rect 1962 95 1966 99
rect 1968 95 1972 99
rect 1974 95 1978 99
rect 1980 95 1984 99
rect 1986 95 1990 99
rect 1962 89 1966 93
rect 1968 89 1972 93
rect 1974 89 1978 93
rect 1980 89 1984 93
rect 1986 89 1990 93
rect 1962 82 1966 86
rect 1968 82 1972 86
rect 1974 82 1978 86
rect 1980 82 1984 86
rect 1986 82 1990 86
rect 1962 76 1966 80
rect 1968 76 1972 80
rect 1974 76 1978 80
rect 1980 76 1984 80
rect 1986 76 1990 80
rect 1962 70 1966 74
rect 1968 70 1972 74
rect 1974 70 1978 74
rect 1980 70 1984 74
rect 1986 70 1990 74
rect 1962 64 1966 68
rect 1968 64 1972 68
rect 1974 64 1978 68
rect 1980 64 1984 68
rect 1986 64 1990 68
rect 2062 95 2066 99
rect 2068 95 2072 99
rect 2074 95 2078 99
rect 2080 95 2084 99
rect 2086 95 2090 99
rect 2062 89 2066 93
rect 2068 89 2072 93
rect 2074 89 2078 93
rect 2080 89 2084 93
rect 2086 89 2090 93
rect 2062 82 2066 86
rect 2068 82 2072 86
rect 2074 82 2078 86
rect 2080 82 2084 86
rect 2086 82 2090 86
rect 2062 76 2066 80
rect 2068 76 2072 80
rect 2074 76 2078 80
rect 2080 76 2084 80
rect 2086 76 2090 80
rect 2062 70 2066 74
rect 2068 70 2072 74
rect 2074 70 2078 74
rect 2080 70 2084 74
rect 2086 70 2090 74
rect 2062 64 2066 68
rect 2068 64 2072 68
rect 2074 64 2078 68
rect 2080 64 2084 68
rect 2086 64 2090 68
rect 1995 53 1999 57
rect 2005 53 2009 57
rect 1961 38 1965 42
rect 1967 38 1971 42
rect 1973 38 1977 42
rect 1979 38 1983 42
rect 1985 38 1989 42
rect 1991 38 1995 42
rect 1997 38 2001 42
rect 1961 20 1965 24
rect 1967 20 1971 24
rect 1973 20 1977 24
rect 1979 20 1983 24
rect 1985 20 1989 24
rect 1991 20 1995 24
rect 1997 20 2001 24
rect 2043 53 2047 57
rect 2053 53 2057 57
rect 2051 38 2055 42
rect 2057 38 2061 42
rect 2063 38 2067 42
rect 2069 38 2073 42
rect 2075 38 2079 42
rect 2081 38 2085 42
rect 2087 38 2091 42
rect 2051 20 2055 24
rect 2057 20 2061 24
rect 2063 20 2067 24
rect 2069 20 2073 24
rect 2075 20 2079 24
rect 2081 20 2085 24
rect 2087 20 2091 24
rect 2435 125 2439 129
rect 2441 125 2445 129
rect 2447 125 2451 129
rect 2453 125 2457 129
rect 2459 125 2463 129
rect 2465 125 2469 129
rect 2471 125 2475 129
rect 2435 112 2439 116
rect 2441 112 2445 116
rect 2447 112 2451 116
rect 2453 112 2457 116
rect 2459 112 2463 116
rect 2465 112 2469 116
rect 2471 112 2475 116
rect 2525 125 2529 129
rect 2531 125 2535 129
rect 2537 125 2541 129
rect 2543 125 2547 129
rect 2549 125 2553 129
rect 2555 125 2559 129
rect 2561 125 2565 129
rect 2525 112 2529 116
rect 2531 112 2535 116
rect 2537 112 2541 116
rect 2543 112 2547 116
rect 2549 112 2553 116
rect 2555 112 2559 116
rect 2561 112 2565 116
rect 2436 95 2440 99
rect 2442 95 2446 99
rect 2448 95 2452 99
rect 2454 95 2458 99
rect 2460 95 2464 99
rect 2436 89 2440 93
rect 2442 89 2446 93
rect 2448 89 2452 93
rect 2454 89 2458 93
rect 2460 89 2464 93
rect 2436 82 2440 86
rect 2442 82 2446 86
rect 2448 82 2452 86
rect 2454 82 2458 86
rect 2460 82 2464 86
rect 2436 76 2440 80
rect 2442 76 2446 80
rect 2448 76 2452 80
rect 2454 76 2458 80
rect 2460 76 2464 80
rect 2436 70 2440 74
rect 2442 70 2446 74
rect 2448 70 2452 74
rect 2454 70 2458 74
rect 2460 70 2464 74
rect 2436 64 2440 68
rect 2442 64 2446 68
rect 2448 64 2452 68
rect 2454 64 2458 68
rect 2460 64 2464 68
rect 2536 95 2540 99
rect 2542 95 2546 99
rect 2548 95 2552 99
rect 2554 95 2558 99
rect 2560 95 2564 99
rect 2536 89 2540 93
rect 2542 89 2546 93
rect 2548 89 2552 93
rect 2554 89 2558 93
rect 2560 89 2564 93
rect 2536 82 2540 86
rect 2542 82 2546 86
rect 2548 82 2552 86
rect 2554 82 2558 86
rect 2560 82 2564 86
rect 2536 76 2540 80
rect 2542 76 2546 80
rect 2548 76 2552 80
rect 2554 76 2558 80
rect 2560 76 2564 80
rect 2536 70 2540 74
rect 2542 70 2546 74
rect 2548 70 2552 74
rect 2554 70 2558 74
rect 2560 70 2564 74
rect 2536 64 2540 68
rect 2542 64 2546 68
rect 2548 64 2552 68
rect 2554 64 2558 68
rect 2560 64 2564 68
rect 2469 53 2473 57
rect 2479 53 2483 57
rect 2435 38 2439 42
rect 2441 38 2445 42
rect 2447 38 2451 42
rect 2453 38 2457 42
rect 2459 38 2463 42
rect 2465 38 2469 42
rect 2471 38 2475 42
rect 2435 20 2439 24
rect 2441 20 2445 24
rect 2447 20 2451 24
rect 2453 20 2457 24
rect 2459 20 2463 24
rect 2465 20 2469 24
rect 2471 20 2475 24
rect 2517 53 2521 57
rect 2527 53 2531 57
rect 2525 38 2529 42
rect 2531 38 2535 42
rect 2537 38 2541 42
rect 2543 38 2547 42
rect 2549 38 2553 42
rect 2555 38 2559 42
rect 2561 38 2565 42
rect 2525 20 2529 24
rect 2531 20 2535 24
rect 2537 20 2541 24
rect 2543 20 2547 24
rect 2549 20 2553 24
rect 2555 20 2559 24
rect 2561 20 2565 24
rect 2909 125 2913 129
rect 2915 125 2919 129
rect 2921 125 2925 129
rect 2927 125 2931 129
rect 2933 125 2937 129
rect 2939 125 2943 129
rect 2945 125 2949 129
rect 2909 112 2913 116
rect 2915 112 2919 116
rect 2921 112 2925 116
rect 2927 112 2931 116
rect 2933 112 2937 116
rect 2939 112 2943 116
rect 2945 112 2949 116
rect 2999 125 3003 129
rect 3005 125 3009 129
rect 3011 125 3015 129
rect 3017 125 3021 129
rect 3023 125 3027 129
rect 3029 125 3033 129
rect 3035 125 3039 129
rect 2999 112 3003 116
rect 3005 112 3009 116
rect 3011 112 3015 116
rect 3017 112 3021 116
rect 3023 112 3027 116
rect 3029 112 3033 116
rect 3035 112 3039 116
rect 2910 95 2914 99
rect 2916 95 2920 99
rect 2922 95 2926 99
rect 2928 95 2932 99
rect 2934 95 2938 99
rect 2910 89 2914 93
rect 2916 89 2920 93
rect 2922 89 2926 93
rect 2928 89 2932 93
rect 2934 89 2938 93
rect 2910 82 2914 86
rect 2916 82 2920 86
rect 2922 82 2926 86
rect 2928 82 2932 86
rect 2934 82 2938 86
rect 2910 76 2914 80
rect 2916 76 2920 80
rect 2922 76 2926 80
rect 2928 76 2932 80
rect 2934 76 2938 80
rect 2910 70 2914 74
rect 2916 70 2920 74
rect 2922 70 2926 74
rect 2928 70 2932 74
rect 2934 70 2938 74
rect 2910 64 2914 68
rect 2916 64 2920 68
rect 2922 64 2926 68
rect 2928 64 2932 68
rect 2934 64 2938 68
rect 3010 95 3014 99
rect 3016 95 3020 99
rect 3022 95 3026 99
rect 3028 95 3032 99
rect 3034 95 3038 99
rect 3010 89 3014 93
rect 3016 89 3020 93
rect 3022 89 3026 93
rect 3028 89 3032 93
rect 3034 89 3038 93
rect 3010 82 3014 86
rect 3016 82 3020 86
rect 3022 82 3026 86
rect 3028 82 3032 86
rect 3034 82 3038 86
rect 3010 76 3014 80
rect 3016 76 3020 80
rect 3022 76 3026 80
rect 3028 76 3032 80
rect 3034 76 3038 80
rect 3010 70 3014 74
rect 3016 70 3020 74
rect 3022 70 3026 74
rect 3028 70 3032 74
rect 3034 70 3038 74
rect 3010 64 3014 68
rect 3016 64 3020 68
rect 3022 64 3026 68
rect 3028 64 3032 68
rect 3034 64 3038 68
rect 2943 53 2947 57
rect 2953 53 2957 57
rect 2909 38 2913 42
rect 2915 38 2919 42
rect 2921 38 2925 42
rect 2927 38 2931 42
rect 2933 38 2937 42
rect 2939 38 2943 42
rect 2945 38 2949 42
rect 2909 20 2913 24
rect 2915 20 2919 24
rect 2921 20 2925 24
rect 2927 20 2931 24
rect 2933 20 2937 24
rect 2939 20 2943 24
rect 2945 20 2949 24
rect 2991 53 2995 57
rect 3001 53 3005 57
rect 2999 38 3003 42
rect 3005 38 3009 42
rect 3011 38 3015 42
rect 3017 38 3021 42
rect 3023 38 3027 42
rect 3029 38 3033 42
rect 3035 38 3039 42
rect 2999 20 3003 24
rect 3005 20 3009 24
rect 3011 20 3015 24
rect 3017 20 3021 24
rect 3023 20 3027 24
rect 3029 20 3033 24
rect 3035 20 3039 24
rect 3383 125 3387 129
rect 3389 125 3393 129
rect 3395 125 3399 129
rect 3401 125 3405 129
rect 3407 125 3411 129
rect 3413 125 3417 129
rect 3419 125 3423 129
rect 3383 112 3387 116
rect 3389 112 3393 116
rect 3395 112 3399 116
rect 3401 112 3405 116
rect 3407 112 3411 116
rect 3413 112 3417 116
rect 3419 112 3423 116
rect 3473 125 3477 129
rect 3479 125 3483 129
rect 3485 125 3489 129
rect 3491 125 3495 129
rect 3497 125 3501 129
rect 3503 125 3507 129
rect 3509 125 3513 129
rect 3473 112 3477 116
rect 3479 112 3483 116
rect 3485 112 3489 116
rect 3491 112 3495 116
rect 3497 112 3501 116
rect 3503 112 3507 116
rect 3509 112 3513 116
rect 3384 95 3388 99
rect 3390 95 3394 99
rect 3396 95 3400 99
rect 3402 95 3406 99
rect 3408 95 3412 99
rect 3384 89 3388 93
rect 3390 89 3394 93
rect 3396 89 3400 93
rect 3402 89 3406 93
rect 3408 89 3412 93
rect 3384 82 3388 86
rect 3390 82 3394 86
rect 3396 82 3400 86
rect 3402 82 3406 86
rect 3408 82 3412 86
rect 3384 76 3388 80
rect 3390 76 3394 80
rect 3396 76 3400 80
rect 3402 76 3406 80
rect 3408 76 3412 80
rect 3384 70 3388 74
rect 3390 70 3394 74
rect 3396 70 3400 74
rect 3402 70 3406 74
rect 3408 70 3412 74
rect 3384 64 3388 68
rect 3390 64 3394 68
rect 3396 64 3400 68
rect 3402 64 3406 68
rect 3408 64 3412 68
rect 3484 95 3488 99
rect 3490 95 3494 99
rect 3496 95 3500 99
rect 3502 95 3506 99
rect 3508 95 3512 99
rect 3484 89 3488 93
rect 3490 89 3494 93
rect 3496 89 3500 93
rect 3502 89 3506 93
rect 3508 89 3512 93
rect 3484 82 3488 86
rect 3490 82 3494 86
rect 3496 82 3500 86
rect 3502 82 3506 86
rect 3508 82 3512 86
rect 3484 76 3488 80
rect 3490 76 3494 80
rect 3496 76 3500 80
rect 3502 76 3506 80
rect 3508 76 3512 80
rect 3484 70 3488 74
rect 3490 70 3494 74
rect 3496 70 3500 74
rect 3502 70 3506 74
rect 3508 70 3512 74
rect 3484 64 3488 68
rect 3490 64 3494 68
rect 3496 64 3500 68
rect 3502 64 3506 68
rect 3508 64 3512 68
rect 3417 53 3421 57
rect 3427 53 3431 57
rect 3383 38 3387 42
rect 3389 38 3393 42
rect 3395 38 3399 42
rect 3401 38 3405 42
rect 3407 38 3411 42
rect 3413 38 3417 42
rect 3419 38 3423 42
rect 3383 20 3387 24
rect 3389 20 3393 24
rect 3395 20 3399 24
rect 3401 20 3405 24
rect 3407 20 3411 24
rect 3413 20 3417 24
rect 3419 20 3423 24
rect 3465 53 3469 57
rect 3475 53 3479 57
rect 3473 38 3477 42
rect 3479 38 3483 42
rect 3485 38 3489 42
rect 3491 38 3495 42
rect 3497 38 3501 42
rect 3503 38 3507 42
rect 3509 38 3513 42
rect 3473 20 3477 24
rect 3479 20 3483 24
rect 3485 20 3489 24
rect 3491 20 3495 24
rect 3497 20 3501 24
rect 3503 20 3507 24
rect 3509 20 3513 24
rect 3857 125 3861 129
rect 3863 125 3867 129
rect 3869 125 3873 129
rect 3875 125 3879 129
rect 3881 125 3885 129
rect 3887 125 3891 129
rect 3893 125 3897 129
rect 3857 112 3861 116
rect 3863 112 3867 116
rect 3869 112 3873 116
rect 3875 112 3879 116
rect 3881 112 3885 116
rect 3887 112 3891 116
rect 3893 112 3897 116
rect 3947 125 3951 129
rect 3953 125 3957 129
rect 3959 125 3963 129
rect 3965 125 3969 129
rect 3971 125 3975 129
rect 3977 125 3981 129
rect 3983 125 3987 129
rect 3947 112 3951 116
rect 3953 112 3957 116
rect 3959 112 3963 116
rect 3965 112 3969 116
rect 3971 112 3975 116
rect 3977 112 3981 116
rect 3983 112 3987 116
rect 3858 95 3862 99
rect 3864 95 3868 99
rect 3870 95 3874 99
rect 3876 95 3880 99
rect 3882 95 3886 99
rect 3858 89 3862 93
rect 3864 89 3868 93
rect 3870 89 3874 93
rect 3876 89 3880 93
rect 3882 89 3886 93
rect 3858 82 3862 86
rect 3864 82 3868 86
rect 3870 82 3874 86
rect 3876 82 3880 86
rect 3882 82 3886 86
rect 3858 76 3862 80
rect 3864 76 3868 80
rect 3870 76 3874 80
rect 3876 76 3880 80
rect 3882 76 3886 80
rect 3858 70 3862 74
rect 3864 70 3868 74
rect 3870 70 3874 74
rect 3876 70 3880 74
rect 3882 70 3886 74
rect 3858 64 3862 68
rect 3864 64 3868 68
rect 3870 64 3874 68
rect 3876 64 3880 68
rect 3882 64 3886 68
rect 3958 95 3962 99
rect 3964 95 3968 99
rect 3970 95 3974 99
rect 3976 95 3980 99
rect 3982 95 3986 99
rect 3958 89 3962 93
rect 3964 89 3968 93
rect 3970 89 3974 93
rect 3976 89 3980 93
rect 3982 89 3986 93
rect 3958 82 3962 86
rect 3964 82 3968 86
rect 3970 82 3974 86
rect 3976 82 3980 86
rect 3982 82 3986 86
rect 3958 76 3962 80
rect 3964 76 3968 80
rect 3970 76 3974 80
rect 3976 76 3980 80
rect 3982 76 3986 80
rect 3958 70 3962 74
rect 3964 70 3968 74
rect 3970 70 3974 74
rect 3976 70 3980 74
rect 3982 70 3986 74
rect 3958 64 3962 68
rect 3964 64 3968 68
rect 3970 64 3974 68
rect 3976 64 3980 68
rect 3982 64 3986 68
rect 3891 53 3895 57
rect 3901 53 3905 57
rect 3857 38 3861 42
rect 3863 38 3867 42
rect 3869 38 3873 42
rect 3875 38 3879 42
rect 3881 38 3885 42
rect 3887 38 3891 42
rect 3893 38 3897 42
rect 3857 20 3861 24
rect 3863 20 3867 24
rect 3869 20 3873 24
rect 3875 20 3879 24
rect 3881 20 3885 24
rect 3887 20 3891 24
rect 3893 20 3897 24
rect 3939 53 3943 57
rect 3949 53 3953 57
rect 3947 38 3951 42
rect 3953 38 3957 42
rect 3959 38 3963 42
rect 3965 38 3969 42
rect 3971 38 3975 42
rect 3977 38 3981 42
rect 3983 38 3987 42
rect 3947 20 3951 24
rect 3953 20 3957 24
rect 3959 20 3963 24
rect 3965 20 3969 24
rect 3971 20 3975 24
rect 3977 20 3981 24
rect 3983 20 3987 24
rect 4331 125 4335 129
rect 4337 125 4341 129
rect 4343 125 4347 129
rect 4349 125 4353 129
rect 4355 125 4359 129
rect 4361 125 4365 129
rect 4367 125 4371 129
rect 4331 112 4335 116
rect 4337 112 4341 116
rect 4343 112 4347 116
rect 4349 112 4353 116
rect 4355 112 4359 116
rect 4361 112 4365 116
rect 4367 112 4371 116
rect 4421 125 4425 129
rect 4427 125 4431 129
rect 4433 125 4437 129
rect 4439 125 4443 129
rect 4445 125 4449 129
rect 4451 125 4455 129
rect 4457 125 4461 129
rect 4421 112 4425 116
rect 4427 112 4431 116
rect 4433 112 4437 116
rect 4439 112 4443 116
rect 4445 112 4449 116
rect 4451 112 4455 116
rect 4457 112 4461 116
rect 4332 95 4336 99
rect 4338 95 4342 99
rect 4344 95 4348 99
rect 4350 95 4354 99
rect 4356 95 4360 99
rect 4332 89 4336 93
rect 4338 89 4342 93
rect 4344 89 4348 93
rect 4350 89 4354 93
rect 4356 89 4360 93
rect 4332 82 4336 86
rect 4338 82 4342 86
rect 4344 82 4348 86
rect 4350 82 4354 86
rect 4356 82 4360 86
rect 4332 76 4336 80
rect 4338 76 4342 80
rect 4344 76 4348 80
rect 4350 76 4354 80
rect 4356 76 4360 80
rect 4332 70 4336 74
rect 4338 70 4342 74
rect 4344 70 4348 74
rect 4350 70 4354 74
rect 4356 70 4360 74
rect 4332 64 4336 68
rect 4338 64 4342 68
rect 4344 64 4348 68
rect 4350 64 4354 68
rect 4356 64 4360 68
rect 4432 95 4436 99
rect 4438 95 4442 99
rect 4444 95 4448 99
rect 4450 95 4454 99
rect 4456 95 4460 99
rect 4432 89 4436 93
rect 4438 89 4442 93
rect 4444 89 4448 93
rect 4450 89 4454 93
rect 4456 89 4460 93
rect 4432 82 4436 86
rect 4438 82 4442 86
rect 4444 82 4448 86
rect 4450 82 4454 86
rect 4456 82 4460 86
rect 4432 76 4436 80
rect 4438 76 4442 80
rect 4444 76 4448 80
rect 4450 76 4454 80
rect 4456 76 4460 80
rect 4432 70 4436 74
rect 4438 70 4442 74
rect 4444 70 4448 74
rect 4450 70 4454 74
rect 4456 70 4460 74
rect 4432 64 4436 68
rect 4438 64 4442 68
rect 4444 64 4448 68
rect 4450 64 4454 68
rect 4456 64 4460 68
rect 4365 53 4369 57
rect 4375 53 4379 57
rect 4331 38 4335 42
rect 4337 38 4341 42
rect 4343 38 4347 42
rect 4349 38 4353 42
rect 4355 38 4359 42
rect 4361 38 4365 42
rect 4367 38 4371 42
rect 4331 20 4335 24
rect 4337 20 4341 24
rect 4343 20 4347 24
rect 4349 20 4353 24
rect 4355 20 4359 24
rect 4361 20 4365 24
rect 4367 20 4371 24
rect 4413 53 4417 57
rect 4423 53 4427 57
rect 4421 38 4425 42
rect 4427 38 4431 42
rect 4433 38 4437 42
rect 4439 38 4443 42
rect 4445 38 4449 42
rect 4451 38 4455 42
rect 4457 38 4461 42
rect 4421 20 4425 24
rect 4427 20 4431 24
rect 4433 20 4437 24
rect 4439 20 4443 24
rect 4445 20 4449 24
rect 4451 20 4455 24
rect 4457 20 4461 24
<< electrodecap >>
rect 376 132 490 137
rect 540 132 668 137
rect 718 132 964 137
rect 1014 132 1142 137
rect 1192 132 1438 137
rect 1488 132 1616 137
rect 1666 132 1912 137
rect 1962 132 2090 137
rect 2140 132 2386 137
rect 2436 132 2564 137
rect 2614 132 2860 137
rect 2910 132 3038 137
rect 3088 132 3334 137
rect 3384 132 3512 137
rect 3562 132 3808 137
rect 3858 132 3986 137
rect 4036 132 4282 137
rect 4332 132 4460 137
rect 4510 132 4624 137
rect 376 105 4624 132
rect 411 62 4589 102
rect 454 51 4546 59
rect 465 17 4535 48
rect 465 12 668 17
rect 718 12 964 17
rect 1014 12 1142 17
rect 1192 12 1438 17
rect 1488 12 1616 17
rect 1666 12 1912 17
rect 1962 12 2090 17
rect 2140 12 2386 17
rect 2436 12 2564 17
rect 2614 12 2860 17
rect 2910 12 3038 17
rect 3088 12 3334 17
rect 3384 12 3512 17
rect 3562 12 3808 17
rect 3858 12 3986 17
rect 4036 12 4282 17
rect 4332 12 4535 17
<< ndiffusion >>
rect 4752 188 4764 189
rect 4752 184 4753 188
rect 4757 184 4759 188
rect 4763 184 4764 188
rect 4752 182 4764 184
rect 4752 178 4753 182
rect 4757 178 4759 182
rect 4763 178 4764 182
rect 4752 176 4764 178
rect 4752 172 4753 176
rect 4757 172 4759 176
rect 4763 172 4764 176
rect 4752 170 4764 172
rect 4752 166 4753 170
rect 4757 166 4759 170
rect 4763 166 4764 170
rect 4752 164 4764 166
rect 4752 160 4753 164
rect 4757 160 4759 164
rect 4763 160 4764 164
rect 4752 158 4764 160
rect 4752 154 4753 158
rect 4757 154 4759 158
rect 4763 154 4764 158
rect 4752 153 4764 154
rect 4778 188 4790 189
rect 4778 184 4779 188
rect 4783 184 4785 188
rect 4789 184 4790 188
rect 4778 182 4790 184
rect 4778 178 4779 182
rect 4783 178 4785 182
rect 4789 178 4790 182
rect 4778 176 4790 178
rect 4778 172 4779 176
rect 4783 172 4785 176
rect 4789 172 4790 176
rect 4778 170 4790 172
rect 4778 166 4779 170
rect 4783 166 4785 170
rect 4789 166 4790 170
rect 4778 164 4790 166
rect 4778 160 4779 164
rect 4783 160 4785 164
rect 4789 160 4790 164
rect 4778 158 4790 160
rect 4778 154 4779 158
rect 4783 154 4785 158
rect 4789 154 4790 158
rect 4778 153 4790 154
<< pdiffusion >>
rect 4652 176 4670 177
rect 4652 172 4653 176
rect 4657 172 4659 176
rect 4663 172 4665 176
rect 4669 172 4670 176
rect 4652 170 4670 172
rect 4652 166 4653 170
rect 4657 166 4659 170
rect 4663 166 4665 170
rect 4669 166 4670 170
rect 4652 165 4670 166
rect 4708 176 4726 177
rect 4708 172 4709 176
rect 4713 172 4715 176
rect 4719 172 4721 176
rect 4725 172 4726 176
rect 4708 170 4726 172
rect 4708 166 4709 170
rect 4713 166 4715 170
rect 4719 166 4721 170
rect 4725 166 4726 170
rect 4708 165 4726 166
<< ndcontact >>
rect 4753 184 4757 188
rect 4759 184 4763 188
rect 4753 178 4757 182
rect 4759 178 4763 182
rect 4753 172 4757 176
rect 4759 172 4763 176
rect 4753 166 4757 170
rect 4759 166 4763 170
rect 4753 160 4757 164
rect 4759 160 4763 164
rect 4753 154 4757 158
rect 4759 154 4763 158
rect 4779 184 4783 188
rect 4785 184 4789 188
rect 4779 178 4783 182
rect 4785 178 4789 182
rect 4779 172 4783 176
rect 4785 172 4789 176
rect 4779 166 4783 170
rect 4785 166 4789 170
rect 4779 160 4783 164
rect 4785 160 4789 164
rect 4779 154 4783 158
rect 4785 154 4789 158
<< pdcontact >>
rect 4653 172 4657 176
rect 4659 172 4663 176
rect 4665 172 4669 176
rect 4653 166 4657 170
rect 4659 166 4663 170
rect 4665 166 4669 170
rect 4709 172 4713 176
rect 4715 172 4719 176
rect 4721 172 4725 176
rect 4709 166 4713 170
rect 4715 166 4719 170
rect 4721 166 4725 170
<< psubstratepdiff >>
rect 364 508 370 511
rect 364 504 365 508
rect 369 504 370 508
rect 364 502 370 504
rect 364 498 365 502
rect 369 498 370 502
rect 364 496 370 498
rect 364 492 365 496
rect 369 492 370 496
rect 364 490 370 492
rect 364 486 365 490
rect 369 486 370 490
rect 364 484 370 486
rect 364 480 365 484
rect 369 480 370 484
rect 364 478 370 480
rect 364 474 365 478
rect 369 474 370 478
rect 364 472 370 474
rect 364 468 365 472
rect 369 468 370 472
rect 364 466 370 468
rect 364 462 365 466
rect 369 462 370 466
rect 364 460 370 462
rect 364 456 365 460
rect 369 456 370 460
rect 364 454 370 456
rect 364 450 365 454
rect 369 450 370 454
rect 364 448 370 450
rect 364 444 365 448
rect 369 444 370 448
rect 364 442 370 444
rect 364 438 365 442
rect 369 438 370 442
rect 364 436 370 438
rect 364 432 365 436
rect 369 432 370 436
rect 364 430 370 432
rect 364 426 365 430
rect 369 426 370 430
rect 364 424 370 426
rect 364 420 365 424
rect 369 420 370 424
rect 364 418 370 420
rect 364 414 365 418
rect 369 414 370 418
rect 364 412 370 414
rect 364 408 365 412
rect 369 408 370 412
rect 364 406 370 408
rect 364 402 365 406
rect 369 402 370 406
rect 364 400 370 402
rect 364 396 365 400
rect 369 396 370 400
rect 364 394 370 396
rect 364 390 365 394
rect 369 390 370 394
rect 364 388 370 390
rect 364 384 365 388
rect 369 384 370 388
rect 364 382 370 384
rect 364 378 365 382
rect 369 378 370 382
rect 364 376 370 378
rect 364 372 365 376
rect 369 372 370 376
rect 364 370 370 372
rect 364 366 365 370
rect 369 366 370 370
rect 364 364 370 366
rect 364 360 365 364
rect 369 360 370 364
rect 364 358 370 360
rect 364 354 365 358
rect 369 354 370 358
rect 364 352 370 354
rect 364 348 365 352
rect 369 348 370 352
rect 364 346 370 348
rect 364 342 365 346
rect 369 342 370 346
rect 364 340 370 342
rect 364 336 365 340
rect 369 336 370 340
rect 364 334 370 336
rect 364 330 365 334
rect 369 330 370 334
rect 364 328 370 330
rect 364 324 365 328
rect 369 324 370 328
rect 364 322 370 324
rect 364 318 365 322
rect 369 318 370 322
rect 364 316 370 318
rect 364 312 365 316
rect 369 312 370 316
rect 364 310 370 312
rect 364 306 365 310
rect 369 306 370 310
rect 364 304 370 306
rect 364 300 365 304
rect 369 300 370 304
rect 364 298 370 300
rect 364 294 365 298
rect 369 294 370 298
rect 364 292 370 294
rect 364 288 365 292
rect 369 288 370 292
rect 364 286 370 288
rect 364 282 365 286
rect 369 282 370 286
rect 364 280 370 282
rect 364 276 365 280
rect 369 276 370 280
rect 364 274 370 276
rect 364 270 365 274
rect 369 270 370 274
rect 364 268 370 270
rect 364 264 365 268
rect 369 264 370 268
rect 364 262 370 264
rect 364 258 365 262
rect 369 258 370 262
rect 364 256 370 258
rect 364 252 365 256
rect 369 252 370 256
rect 364 250 370 252
rect 364 246 365 250
rect 369 246 370 250
rect 364 244 370 246
rect 364 240 365 244
rect 369 240 370 244
rect 364 238 370 240
rect 364 234 365 238
rect 369 234 370 238
rect 364 232 370 234
rect 364 228 365 232
rect 369 228 370 232
rect 364 226 370 228
rect 364 222 365 226
rect 369 222 370 226
rect 364 220 370 222
rect 364 216 365 220
rect 369 216 370 220
rect 364 214 370 216
rect 364 210 365 214
rect 369 210 370 214
rect 364 208 370 210
rect 364 204 365 208
rect 369 204 370 208
rect 364 202 370 204
rect 364 198 365 202
rect 369 198 370 202
rect 364 196 370 198
rect 364 192 365 196
rect 369 192 370 196
rect 364 190 370 192
rect 364 186 365 190
rect 369 186 370 190
rect 364 184 370 186
rect 364 180 365 184
rect 369 180 370 184
rect 364 178 370 180
rect 364 174 365 178
rect 369 174 370 178
rect 364 172 370 174
rect 364 168 365 172
rect 369 168 370 172
rect 364 166 370 168
rect 364 162 365 166
rect 369 162 370 166
rect 364 160 370 162
rect 364 156 365 160
rect 369 156 370 160
rect 364 154 370 156
rect 364 150 365 154
rect 369 150 370 154
rect 364 149 370 150
rect 838 508 844 511
rect 838 504 839 508
rect 843 504 844 508
rect 838 502 844 504
rect 838 498 839 502
rect 843 498 844 502
rect 838 496 844 498
rect 838 492 839 496
rect 843 492 844 496
rect 838 490 844 492
rect 838 486 839 490
rect 843 486 844 490
rect 838 484 844 486
rect 838 480 839 484
rect 843 480 844 484
rect 838 478 844 480
rect 838 474 839 478
rect 843 474 844 478
rect 838 472 844 474
rect 838 468 839 472
rect 843 468 844 472
rect 838 466 844 468
rect 838 462 839 466
rect 843 462 844 466
rect 838 460 844 462
rect 838 456 839 460
rect 843 456 844 460
rect 838 454 844 456
rect 838 450 839 454
rect 843 450 844 454
rect 838 448 844 450
rect 838 444 839 448
rect 843 444 844 448
rect 838 442 844 444
rect 838 438 839 442
rect 843 438 844 442
rect 838 436 844 438
rect 838 432 839 436
rect 843 432 844 436
rect 838 430 844 432
rect 838 426 839 430
rect 843 426 844 430
rect 838 424 844 426
rect 838 420 839 424
rect 843 420 844 424
rect 838 418 844 420
rect 838 414 839 418
rect 843 414 844 418
rect 838 412 844 414
rect 838 408 839 412
rect 843 408 844 412
rect 838 406 844 408
rect 838 402 839 406
rect 843 402 844 406
rect 838 400 844 402
rect 838 396 839 400
rect 843 396 844 400
rect 838 394 844 396
rect 838 390 839 394
rect 843 390 844 394
rect 838 388 844 390
rect 838 384 839 388
rect 843 384 844 388
rect 838 382 844 384
rect 838 378 839 382
rect 843 378 844 382
rect 838 376 844 378
rect 838 372 839 376
rect 843 372 844 376
rect 838 370 844 372
rect 838 366 839 370
rect 843 366 844 370
rect 838 364 844 366
rect 838 360 839 364
rect 843 360 844 364
rect 838 358 844 360
rect 838 354 839 358
rect 843 354 844 358
rect 838 352 844 354
rect 838 348 839 352
rect 843 348 844 352
rect 838 346 844 348
rect 838 342 839 346
rect 843 342 844 346
rect 838 340 844 342
rect 838 336 839 340
rect 843 336 844 340
rect 838 334 844 336
rect 838 330 839 334
rect 843 330 844 334
rect 838 328 844 330
rect 838 324 839 328
rect 843 324 844 328
rect 838 322 844 324
rect 838 318 839 322
rect 843 318 844 322
rect 838 316 844 318
rect 838 312 839 316
rect 843 312 844 316
rect 838 310 844 312
rect 838 306 839 310
rect 843 306 844 310
rect 838 304 844 306
rect 838 300 839 304
rect 843 300 844 304
rect 838 298 844 300
rect 838 294 839 298
rect 843 294 844 298
rect 838 292 844 294
rect 838 288 839 292
rect 843 288 844 292
rect 838 286 844 288
rect 838 282 839 286
rect 843 282 844 286
rect 838 280 844 282
rect 838 276 839 280
rect 843 276 844 280
rect 838 274 844 276
rect 838 270 839 274
rect 843 270 844 274
rect 838 268 844 270
rect 838 264 839 268
rect 843 264 844 268
rect 838 262 844 264
rect 838 258 839 262
rect 843 258 844 262
rect 838 256 844 258
rect 838 252 839 256
rect 843 252 844 256
rect 838 250 844 252
rect 838 246 839 250
rect 843 246 844 250
rect 838 244 844 246
rect 838 240 839 244
rect 843 240 844 244
rect 838 238 844 240
rect 838 234 839 238
rect 843 234 844 238
rect 838 232 844 234
rect 838 228 839 232
rect 843 228 844 232
rect 838 226 844 228
rect 838 222 839 226
rect 843 222 844 226
rect 838 220 844 222
rect 838 216 839 220
rect 843 216 844 220
rect 838 214 844 216
rect 838 210 839 214
rect 843 210 844 214
rect 838 208 844 210
rect 838 204 839 208
rect 843 204 844 208
rect 838 202 844 204
rect 838 198 839 202
rect 843 198 844 202
rect 838 196 844 198
rect 838 192 839 196
rect 843 192 844 196
rect 838 190 844 192
rect 838 186 839 190
rect 843 186 844 190
rect 838 184 844 186
rect 838 180 839 184
rect 843 180 844 184
rect 838 178 844 180
rect 838 174 839 178
rect 843 174 844 178
rect 838 172 844 174
rect 838 168 839 172
rect 843 168 844 172
rect 838 166 844 168
rect 838 162 839 166
rect 843 162 844 166
rect 838 160 844 162
rect 838 156 839 160
rect 843 156 844 160
rect 838 154 844 156
rect 838 150 839 154
rect 843 150 844 154
rect 838 149 844 150
rect 1312 508 1318 511
rect 1312 504 1313 508
rect 1317 504 1318 508
rect 1312 502 1318 504
rect 1312 498 1313 502
rect 1317 498 1318 502
rect 1312 496 1318 498
rect 1312 492 1313 496
rect 1317 492 1318 496
rect 1312 490 1318 492
rect 1312 486 1313 490
rect 1317 486 1318 490
rect 1312 484 1318 486
rect 1312 480 1313 484
rect 1317 480 1318 484
rect 1312 478 1318 480
rect 1312 474 1313 478
rect 1317 474 1318 478
rect 1312 472 1318 474
rect 1312 468 1313 472
rect 1317 468 1318 472
rect 1312 466 1318 468
rect 1312 462 1313 466
rect 1317 462 1318 466
rect 1312 460 1318 462
rect 1312 456 1313 460
rect 1317 456 1318 460
rect 1312 454 1318 456
rect 1312 450 1313 454
rect 1317 450 1318 454
rect 1312 448 1318 450
rect 1312 444 1313 448
rect 1317 444 1318 448
rect 1312 442 1318 444
rect 1312 438 1313 442
rect 1317 438 1318 442
rect 1312 436 1318 438
rect 1312 432 1313 436
rect 1317 432 1318 436
rect 1312 430 1318 432
rect 1312 426 1313 430
rect 1317 426 1318 430
rect 1312 424 1318 426
rect 1312 420 1313 424
rect 1317 420 1318 424
rect 1312 418 1318 420
rect 1312 414 1313 418
rect 1317 414 1318 418
rect 1312 412 1318 414
rect 1312 408 1313 412
rect 1317 408 1318 412
rect 1312 406 1318 408
rect 1312 402 1313 406
rect 1317 402 1318 406
rect 1312 400 1318 402
rect 1312 396 1313 400
rect 1317 396 1318 400
rect 1312 394 1318 396
rect 1312 390 1313 394
rect 1317 390 1318 394
rect 1312 388 1318 390
rect 1312 384 1313 388
rect 1317 384 1318 388
rect 1312 382 1318 384
rect 1312 378 1313 382
rect 1317 378 1318 382
rect 1312 376 1318 378
rect 1312 372 1313 376
rect 1317 372 1318 376
rect 1312 370 1318 372
rect 1312 366 1313 370
rect 1317 366 1318 370
rect 1312 364 1318 366
rect 1312 360 1313 364
rect 1317 360 1318 364
rect 1312 358 1318 360
rect 1312 354 1313 358
rect 1317 354 1318 358
rect 1312 352 1318 354
rect 1312 348 1313 352
rect 1317 348 1318 352
rect 1312 346 1318 348
rect 1312 342 1313 346
rect 1317 342 1318 346
rect 1312 340 1318 342
rect 1312 336 1313 340
rect 1317 336 1318 340
rect 1312 334 1318 336
rect 1312 330 1313 334
rect 1317 330 1318 334
rect 1312 328 1318 330
rect 1312 324 1313 328
rect 1317 324 1318 328
rect 1312 322 1318 324
rect 1312 318 1313 322
rect 1317 318 1318 322
rect 1312 316 1318 318
rect 1312 312 1313 316
rect 1317 312 1318 316
rect 1312 310 1318 312
rect 1312 306 1313 310
rect 1317 306 1318 310
rect 1312 304 1318 306
rect 1312 300 1313 304
rect 1317 300 1318 304
rect 1312 298 1318 300
rect 1312 294 1313 298
rect 1317 294 1318 298
rect 1312 292 1318 294
rect 1312 288 1313 292
rect 1317 288 1318 292
rect 1312 286 1318 288
rect 1312 282 1313 286
rect 1317 282 1318 286
rect 1312 280 1318 282
rect 1312 276 1313 280
rect 1317 276 1318 280
rect 1312 274 1318 276
rect 1312 270 1313 274
rect 1317 270 1318 274
rect 1312 268 1318 270
rect 1312 264 1313 268
rect 1317 264 1318 268
rect 1312 262 1318 264
rect 1312 258 1313 262
rect 1317 258 1318 262
rect 1312 256 1318 258
rect 1312 252 1313 256
rect 1317 252 1318 256
rect 1312 250 1318 252
rect 1312 246 1313 250
rect 1317 246 1318 250
rect 1312 244 1318 246
rect 1312 240 1313 244
rect 1317 240 1318 244
rect 1312 238 1318 240
rect 1312 234 1313 238
rect 1317 234 1318 238
rect 1312 232 1318 234
rect 1312 228 1313 232
rect 1317 228 1318 232
rect 1312 226 1318 228
rect 1312 222 1313 226
rect 1317 222 1318 226
rect 1312 220 1318 222
rect 1312 216 1313 220
rect 1317 216 1318 220
rect 1312 214 1318 216
rect 1312 210 1313 214
rect 1317 210 1318 214
rect 1312 208 1318 210
rect 1312 204 1313 208
rect 1317 204 1318 208
rect 1312 202 1318 204
rect 1312 198 1313 202
rect 1317 198 1318 202
rect 1312 196 1318 198
rect 1312 192 1313 196
rect 1317 192 1318 196
rect 1312 190 1318 192
rect 1312 186 1313 190
rect 1317 186 1318 190
rect 1312 184 1318 186
rect 1312 180 1313 184
rect 1317 180 1318 184
rect 1312 178 1318 180
rect 1312 174 1313 178
rect 1317 174 1318 178
rect 1312 172 1318 174
rect 1312 168 1313 172
rect 1317 168 1318 172
rect 1312 166 1318 168
rect 1312 162 1313 166
rect 1317 162 1318 166
rect 1312 160 1318 162
rect 1312 156 1313 160
rect 1317 156 1318 160
rect 1312 154 1318 156
rect 1312 150 1313 154
rect 1317 150 1318 154
rect 1312 149 1318 150
rect 1786 508 1792 511
rect 1786 504 1787 508
rect 1791 504 1792 508
rect 1786 502 1792 504
rect 1786 498 1787 502
rect 1791 498 1792 502
rect 1786 496 1792 498
rect 1786 492 1787 496
rect 1791 492 1792 496
rect 1786 490 1792 492
rect 1786 486 1787 490
rect 1791 486 1792 490
rect 1786 484 1792 486
rect 1786 480 1787 484
rect 1791 480 1792 484
rect 1786 478 1792 480
rect 1786 474 1787 478
rect 1791 474 1792 478
rect 1786 472 1792 474
rect 1786 468 1787 472
rect 1791 468 1792 472
rect 1786 466 1792 468
rect 1786 462 1787 466
rect 1791 462 1792 466
rect 1786 460 1792 462
rect 1786 456 1787 460
rect 1791 456 1792 460
rect 1786 454 1792 456
rect 1786 450 1787 454
rect 1791 450 1792 454
rect 1786 448 1792 450
rect 1786 444 1787 448
rect 1791 444 1792 448
rect 1786 442 1792 444
rect 1786 438 1787 442
rect 1791 438 1792 442
rect 1786 436 1792 438
rect 1786 432 1787 436
rect 1791 432 1792 436
rect 1786 430 1792 432
rect 1786 426 1787 430
rect 1791 426 1792 430
rect 1786 424 1792 426
rect 1786 420 1787 424
rect 1791 420 1792 424
rect 1786 418 1792 420
rect 1786 414 1787 418
rect 1791 414 1792 418
rect 1786 412 1792 414
rect 1786 408 1787 412
rect 1791 408 1792 412
rect 1786 406 1792 408
rect 1786 402 1787 406
rect 1791 402 1792 406
rect 1786 400 1792 402
rect 1786 396 1787 400
rect 1791 396 1792 400
rect 1786 394 1792 396
rect 1786 390 1787 394
rect 1791 390 1792 394
rect 1786 388 1792 390
rect 1786 384 1787 388
rect 1791 384 1792 388
rect 1786 382 1792 384
rect 1786 378 1787 382
rect 1791 378 1792 382
rect 1786 376 1792 378
rect 1786 372 1787 376
rect 1791 372 1792 376
rect 1786 370 1792 372
rect 1786 366 1787 370
rect 1791 366 1792 370
rect 1786 364 1792 366
rect 1786 360 1787 364
rect 1791 360 1792 364
rect 1786 358 1792 360
rect 1786 354 1787 358
rect 1791 354 1792 358
rect 1786 352 1792 354
rect 1786 348 1787 352
rect 1791 348 1792 352
rect 1786 346 1792 348
rect 1786 342 1787 346
rect 1791 342 1792 346
rect 1786 340 1792 342
rect 1786 336 1787 340
rect 1791 336 1792 340
rect 1786 334 1792 336
rect 1786 330 1787 334
rect 1791 330 1792 334
rect 1786 328 1792 330
rect 1786 324 1787 328
rect 1791 324 1792 328
rect 1786 322 1792 324
rect 1786 318 1787 322
rect 1791 318 1792 322
rect 1786 316 1792 318
rect 1786 312 1787 316
rect 1791 312 1792 316
rect 1786 310 1792 312
rect 1786 306 1787 310
rect 1791 306 1792 310
rect 1786 304 1792 306
rect 1786 300 1787 304
rect 1791 300 1792 304
rect 1786 298 1792 300
rect 1786 294 1787 298
rect 1791 294 1792 298
rect 1786 292 1792 294
rect 1786 288 1787 292
rect 1791 288 1792 292
rect 1786 286 1792 288
rect 1786 282 1787 286
rect 1791 282 1792 286
rect 1786 280 1792 282
rect 1786 276 1787 280
rect 1791 276 1792 280
rect 1786 274 1792 276
rect 1786 270 1787 274
rect 1791 270 1792 274
rect 1786 268 1792 270
rect 1786 264 1787 268
rect 1791 264 1792 268
rect 1786 262 1792 264
rect 1786 258 1787 262
rect 1791 258 1792 262
rect 1786 256 1792 258
rect 1786 252 1787 256
rect 1791 252 1792 256
rect 1786 250 1792 252
rect 1786 246 1787 250
rect 1791 246 1792 250
rect 1786 244 1792 246
rect 1786 240 1787 244
rect 1791 240 1792 244
rect 1786 238 1792 240
rect 1786 234 1787 238
rect 1791 234 1792 238
rect 1786 232 1792 234
rect 1786 228 1787 232
rect 1791 228 1792 232
rect 1786 226 1792 228
rect 1786 222 1787 226
rect 1791 222 1792 226
rect 1786 220 1792 222
rect 1786 216 1787 220
rect 1791 216 1792 220
rect 1786 214 1792 216
rect 1786 210 1787 214
rect 1791 210 1792 214
rect 1786 208 1792 210
rect 1786 204 1787 208
rect 1791 204 1792 208
rect 1786 202 1792 204
rect 1786 198 1787 202
rect 1791 198 1792 202
rect 1786 196 1792 198
rect 1786 192 1787 196
rect 1791 192 1792 196
rect 1786 190 1792 192
rect 1786 186 1787 190
rect 1791 186 1792 190
rect 1786 184 1792 186
rect 1786 180 1787 184
rect 1791 180 1792 184
rect 1786 178 1792 180
rect 1786 174 1787 178
rect 1791 174 1792 178
rect 1786 172 1792 174
rect 1786 168 1787 172
rect 1791 168 1792 172
rect 1786 166 1792 168
rect 1786 162 1787 166
rect 1791 162 1792 166
rect 1786 160 1792 162
rect 1786 156 1787 160
rect 1791 156 1792 160
rect 1786 154 1792 156
rect 1786 150 1787 154
rect 1791 150 1792 154
rect 1786 149 1792 150
rect 2260 508 2266 511
rect 2260 504 2261 508
rect 2265 504 2266 508
rect 2260 502 2266 504
rect 2260 498 2261 502
rect 2265 498 2266 502
rect 2260 496 2266 498
rect 2260 492 2261 496
rect 2265 492 2266 496
rect 2260 490 2266 492
rect 2260 486 2261 490
rect 2265 486 2266 490
rect 2260 484 2266 486
rect 2260 480 2261 484
rect 2265 480 2266 484
rect 2260 478 2266 480
rect 2260 474 2261 478
rect 2265 474 2266 478
rect 2260 472 2266 474
rect 2260 468 2261 472
rect 2265 468 2266 472
rect 2260 466 2266 468
rect 2260 462 2261 466
rect 2265 462 2266 466
rect 2260 460 2266 462
rect 2260 456 2261 460
rect 2265 456 2266 460
rect 2260 454 2266 456
rect 2260 450 2261 454
rect 2265 450 2266 454
rect 2260 448 2266 450
rect 2260 444 2261 448
rect 2265 444 2266 448
rect 2260 442 2266 444
rect 2260 438 2261 442
rect 2265 438 2266 442
rect 2260 436 2266 438
rect 2260 432 2261 436
rect 2265 432 2266 436
rect 2260 430 2266 432
rect 2260 426 2261 430
rect 2265 426 2266 430
rect 2260 424 2266 426
rect 2260 420 2261 424
rect 2265 420 2266 424
rect 2260 418 2266 420
rect 2260 414 2261 418
rect 2265 414 2266 418
rect 2260 412 2266 414
rect 2260 408 2261 412
rect 2265 408 2266 412
rect 2260 406 2266 408
rect 2260 402 2261 406
rect 2265 402 2266 406
rect 2260 400 2266 402
rect 2260 396 2261 400
rect 2265 396 2266 400
rect 2260 394 2266 396
rect 2260 390 2261 394
rect 2265 390 2266 394
rect 2260 388 2266 390
rect 2260 384 2261 388
rect 2265 384 2266 388
rect 2260 382 2266 384
rect 2260 378 2261 382
rect 2265 378 2266 382
rect 2260 376 2266 378
rect 2260 372 2261 376
rect 2265 372 2266 376
rect 2260 370 2266 372
rect 2260 366 2261 370
rect 2265 366 2266 370
rect 2260 364 2266 366
rect 2260 360 2261 364
rect 2265 360 2266 364
rect 2260 358 2266 360
rect 2260 354 2261 358
rect 2265 354 2266 358
rect 2260 352 2266 354
rect 2260 348 2261 352
rect 2265 348 2266 352
rect 2260 346 2266 348
rect 2260 342 2261 346
rect 2265 342 2266 346
rect 2260 340 2266 342
rect 2260 336 2261 340
rect 2265 336 2266 340
rect 2260 334 2266 336
rect 2260 330 2261 334
rect 2265 330 2266 334
rect 2260 328 2266 330
rect 2260 324 2261 328
rect 2265 324 2266 328
rect 2260 322 2266 324
rect 2260 318 2261 322
rect 2265 318 2266 322
rect 2260 316 2266 318
rect 2260 312 2261 316
rect 2265 312 2266 316
rect 2260 310 2266 312
rect 2260 306 2261 310
rect 2265 306 2266 310
rect 2260 304 2266 306
rect 2260 300 2261 304
rect 2265 300 2266 304
rect 2260 298 2266 300
rect 2260 294 2261 298
rect 2265 294 2266 298
rect 2260 292 2266 294
rect 2260 288 2261 292
rect 2265 288 2266 292
rect 2260 286 2266 288
rect 2260 282 2261 286
rect 2265 282 2266 286
rect 2260 280 2266 282
rect 2260 276 2261 280
rect 2265 276 2266 280
rect 2260 274 2266 276
rect 2260 270 2261 274
rect 2265 270 2266 274
rect 2260 268 2266 270
rect 2260 264 2261 268
rect 2265 264 2266 268
rect 2260 262 2266 264
rect 2260 258 2261 262
rect 2265 258 2266 262
rect 2260 256 2266 258
rect 2260 252 2261 256
rect 2265 252 2266 256
rect 2260 250 2266 252
rect 2260 246 2261 250
rect 2265 246 2266 250
rect 2260 244 2266 246
rect 2260 240 2261 244
rect 2265 240 2266 244
rect 2260 238 2266 240
rect 2260 234 2261 238
rect 2265 234 2266 238
rect 2260 232 2266 234
rect 2260 228 2261 232
rect 2265 228 2266 232
rect 2260 226 2266 228
rect 2260 222 2261 226
rect 2265 222 2266 226
rect 2260 220 2266 222
rect 2260 216 2261 220
rect 2265 216 2266 220
rect 2260 214 2266 216
rect 2260 210 2261 214
rect 2265 210 2266 214
rect 2260 208 2266 210
rect 2260 204 2261 208
rect 2265 204 2266 208
rect 2260 202 2266 204
rect 2260 198 2261 202
rect 2265 198 2266 202
rect 2260 196 2266 198
rect 2260 192 2261 196
rect 2265 192 2266 196
rect 2260 190 2266 192
rect 2260 186 2261 190
rect 2265 186 2266 190
rect 2260 184 2266 186
rect 2260 180 2261 184
rect 2265 180 2266 184
rect 2260 178 2266 180
rect 2260 174 2261 178
rect 2265 174 2266 178
rect 2260 172 2266 174
rect 2260 168 2261 172
rect 2265 168 2266 172
rect 2260 166 2266 168
rect 2260 162 2261 166
rect 2265 162 2266 166
rect 2260 160 2266 162
rect 2260 156 2261 160
rect 2265 156 2266 160
rect 2260 154 2266 156
rect 2260 150 2261 154
rect 2265 150 2266 154
rect 2260 149 2266 150
rect 2734 508 2740 511
rect 2734 504 2735 508
rect 2739 504 2740 508
rect 2734 502 2740 504
rect 2734 498 2735 502
rect 2739 498 2740 502
rect 2734 496 2740 498
rect 2734 492 2735 496
rect 2739 492 2740 496
rect 2734 490 2740 492
rect 2734 486 2735 490
rect 2739 486 2740 490
rect 2734 484 2740 486
rect 2734 480 2735 484
rect 2739 480 2740 484
rect 2734 478 2740 480
rect 2734 474 2735 478
rect 2739 474 2740 478
rect 2734 472 2740 474
rect 2734 468 2735 472
rect 2739 468 2740 472
rect 2734 466 2740 468
rect 2734 462 2735 466
rect 2739 462 2740 466
rect 2734 460 2740 462
rect 2734 456 2735 460
rect 2739 456 2740 460
rect 2734 454 2740 456
rect 2734 450 2735 454
rect 2739 450 2740 454
rect 2734 448 2740 450
rect 2734 444 2735 448
rect 2739 444 2740 448
rect 2734 442 2740 444
rect 2734 438 2735 442
rect 2739 438 2740 442
rect 2734 436 2740 438
rect 2734 432 2735 436
rect 2739 432 2740 436
rect 2734 430 2740 432
rect 2734 426 2735 430
rect 2739 426 2740 430
rect 2734 424 2740 426
rect 2734 420 2735 424
rect 2739 420 2740 424
rect 2734 418 2740 420
rect 2734 414 2735 418
rect 2739 414 2740 418
rect 2734 412 2740 414
rect 2734 408 2735 412
rect 2739 408 2740 412
rect 2734 406 2740 408
rect 2734 402 2735 406
rect 2739 402 2740 406
rect 2734 400 2740 402
rect 2734 396 2735 400
rect 2739 396 2740 400
rect 2734 394 2740 396
rect 2734 390 2735 394
rect 2739 390 2740 394
rect 2734 388 2740 390
rect 2734 384 2735 388
rect 2739 384 2740 388
rect 2734 382 2740 384
rect 2734 378 2735 382
rect 2739 378 2740 382
rect 2734 376 2740 378
rect 2734 372 2735 376
rect 2739 372 2740 376
rect 2734 370 2740 372
rect 2734 366 2735 370
rect 2739 366 2740 370
rect 2734 364 2740 366
rect 2734 360 2735 364
rect 2739 360 2740 364
rect 2734 358 2740 360
rect 2734 354 2735 358
rect 2739 354 2740 358
rect 2734 352 2740 354
rect 2734 348 2735 352
rect 2739 348 2740 352
rect 2734 346 2740 348
rect 2734 342 2735 346
rect 2739 342 2740 346
rect 2734 340 2740 342
rect 2734 336 2735 340
rect 2739 336 2740 340
rect 2734 334 2740 336
rect 2734 330 2735 334
rect 2739 330 2740 334
rect 2734 328 2740 330
rect 2734 324 2735 328
rect 2739 324 2740 328
rect 2734 322 2740 324
rect 2734 318 2735 322
rect 2739 318 2740 322
rect 2734 316 2740 318
rect 2734 312 2735 316
rect 2739 312 2740 316
rect 2734 310 2740 312
rect 2734 306 2735 310
rect 2739 306 2740 310
rect 2734 304 2740 306
rect 2734 300 2735 304
rect 2739 300 2740 304
rect 2734 298 2740 300
rect 2734 294 2735 298
rect 2739 294 2740 298
rect 2734 292 2740 294
rect 2734 288 2735 292
rect 2739 288 2740 292
rect 2734 286 2740 288
rect 2734 282 2735 286
rect 2739 282 2740 286
rect 2734 280 2740 282
rect 2734 276 2735 280
rect 2739 276 2740 280
rect 2734 274 2740 276
rect 2734 270 2735 274
rect 2739 270 2740 274
rect 2734 268 2740 270
rect 2734 264 2735 268
rect 2739 264 2740 268
rect 2734 262 2740 264
rect 2734 258 2735 262
rect 2739 258 2740 262
rect 2734 256 2740 258
rect 2734 252 2735 256
rect 2739 252 2740 256
rect 2734 250 2740 252
rect 2734 246 2735 250
rect 2739 246 2740 250
rect 2734 244 2740 246
rect 2734 240 2735 244
rect 2739 240 2740 244
rect 2734 238 2740 240
rect 2734 234 2735 238
rect 2739 234 2740 238
rect 2734 232 2740 234
rect 2734 228 2735 232
rect 2739 228 2740 232
rect 2734 226 2740 228
rect 2734 222 2735 226
rect 2739 222 2740 226
rect 2734 220 2740 222
rect 2734 216 2735 220
rect 2739 216 2740 220
rect 2734 214 2740 216
rect 2734 210 2735 214
rect 2739 210 2740 214
rect 2734 208 2740 210
rect 2734 204 2735 208
rect 2739 204 2740 208
rect 2734 202 2740 204
rect 2734 198 2735 202
rect 2739 198 2740 202
rect 2734 196 2740 198
rect 2734 192 2735 196
rect 2739 192 2740 196
rect 2734 190 2740 192
rect 2734 186 2735 190
rect 2739 186 2740 190
rect 2734 184 2740 186
rect 2734 180 2735 184
rect 2739 180 2740 184
rect 2734 178 2740 180
rect 2734 174 2735 178
rect 2739 174 2740 178
rect 2734 172 2740 174
rect 2734 168 2735 172
rect 2739 168 2740 172
rect 2734 166 2740 168
rect 2734 162 2735 166
rect 2739 162 2740 166
rect 2734 160 2740 162
rect 2734 156 2735 160
rect 2739 156 2740 160
rect 2734 154 2740 156
rect 2734 150 2735 154
rect 2739 150 2740 154
rect 2734 149 2740 150
rect 3208 508 3214 511
rect 3208 504 3209 508
rect 3213 504 3214 508
rect 3208 502 3214 504
rect 3208 498 3209 502
rect 3213 498 3214 502
rect 3208 496 3214 498
rect 3208 492 3209 496
rect 3213 492 3214 496
rect 3208 490 3214 492
rect 3208 486 3209 490
rect 3213 486 3214 490
rect 3208 484 3214 486
rect 3208 480 3209 484
rect 3213 480 3214 484
rect 3208 478 3214 480
rect 3208 474 3209 478
rect 3213 474 3214 478
rect 3208 472 3214 474
rect 3208 468 3209 472
rect 3213 468 3214 472
rect 3208 466 3214 468
rect 3208 462 3209 466
rect 3213 462 3214 466
rect 3208 460 3214 462
rect 3208 456 3209 460
rect 3213 456 3214 460
rect 3208 454 3214 456
rect 3208 450 3209 454
rect 3213 450 3214 454
rect 3208 448 3214 450
rect 3208 444 3209 448
rect 3213 444 3214 448
rect 3208 442 3214 444
rect 3208 438 3209 442
rect 3213 438 3214 442
rect 3208 436 3214 438
rect 3208 432 3209 436
rect 3213 432 3214 436
rect 3208 430 3214 432
rect 3208 426 3209 430
rect 3213 426 3214 430
rect 3208 424 3214 426
rect 3208 420 3209 424
rect 3213 420 3214 424
rect 3208 418 3214 420
rect 3208 414 3209 418
rect 3213 414 3214 418
rect 3208 412 3214 414
rect 3208 408 3209 412
rect 3213 408 3214 412
rect 3208 406 3214 408
rect 3208 402 3209 406
rect 3213 402 3214 406
rect 3208 400 3214 402
rect 3208 396 3209 400
rect 3213 396 3214 400
rect 3208 394 3214 396
rect 3208 390 3209 394
rect 3213 390 3214 394
rect 3208 388 3214 390
rect 3208 384 3209 388
rect 3213 384 3214 388
rect 3208 382 3214 384
rect 3208 378 3209 382
rect 3213 378 3214 382
rect 3208 376 3214 378
rect 3208 372 3209 376
rect 3213 372 3214 376
rect 3208 370 3214 372
rect 3208 366 3209 370
rect 3213 366 3214 370
rect 3208 364 3214 366
rect 3208 360 3209 364
rect 3213 360 3214 364
rect 3208 358 3214 360
rect 3208 354 3209 358
rect 3213 354 3214 358
rect 3208 352 3214 354
rect 3208 348 3209 352
rect 3213 348 3214 352
rect 3208 346 3214 348
rect 3208 342 3209 346
rect 3213 342 3214 346
rect 3208 340 3214 342
rect 3208 336 3209 340
rect 3213 336 3214 340
rect 3208 334 3214 336
rect 3208 330 3209 334
rect 3213 330 3214 334
rect 3208 328 3214 330
rect 3208 324 3209 328
rect 3213 324 3214 328
rect 3208 322 3214 324
rect 3208 318 3209 322
rect 3213 318 3214 322
rect 3208 316 3214 318
rect 3208 312 3209 316
rect 3213 312 3214 316
rect 3208 310 3214 312
rect 3208 306 3209 310
rect 3213 306 3214 310
rect 3208 304 3214 306
rect 3208 300 3209 304
rect 3213 300 3214 304
rect 3208 298 3214 300
rect 3208 294 3209 298
rect 3213 294 3214 298
rect 3208 292 3214 294
rect 3208 288 3209 292
rect 3213 288 3214 292
rect 3208 286 3214 288
rect 3208 282 3209 286
rect 3213 282 3214 286
rect 3208 280 3214 282
rect 3208 276 3209 280
rect 3213 276 3214 280
rect 3208 274 3214 276
rect 3208 270 3209 274
rect 3213 270 3214 274
rect 3208 268 3214 270
rect 3208 264 3209 268
rect 3213 264 3214 268
rect 3208 262 3214 264
rect 3208 258 3209 262
rect 3213 258 3214 262
rect 3208 256 3214 258
rect 3208 252 3209 256
rect 3213 252 3214 256
rect 3208 250 3214 252
rect 3208 246 3209 250
rect 3213 246 3214 250
rect 3208 244 3214 246
rect 3208 240 3209 244
rect 3213 240 3214 244
rect 3208 238 3214 240
rect 3208 234 3209 238
rect 3213 234 3214 238
rect 3208 232 3214 234
rect 3208 228 3209 232
rect 3213 228 3214 232
rect 3208 226 3214 228
rect 3208 222 3209 226
rect 3213 222 3214 226
rect 3208 220 3214 222
rect 3208 216 3209 220
rect 3213 216 3214 220
rect 3208 214 3214 216
rect 3208 210 3209 214
rect 3213 210 3214 214
rect 3208 208 3214 210
rect 3208 204 3209 208
rect 3213 204 3214 208
rect 3208 202 3214 204
rect 3208 198 3209 202
rect 3213 198 3214 202
rect 3208 196 3214 198
rect 3208 192 3209 196
rect 3213 192 3214 196
rect 3208 190 3214 192
rect 3208 186 3209 190
rect 3213 186 3214 190
rect 3208 184 3214 186
rect 3208 180 3209 184
rect 3213 180 3214 184
rect 3208 178 3214 180
rect 3208 174 3209 178
rect 3213 174 3214 178
rect 3208 172 3214 174
rect 3208 168 3209 172
rect 3213 168 3214 172
rect 3208 166 3214 168
rect 3208 162 3209 166
rect 3213 162 3214 166
rect 3208 160 3214 162
rect 3208 156 3209 160
rect 3213 156 3214 160
rect 3208 154 3214 156
rect 3208 150 3209 154
rect 3213 150 3214 154
rect 3208 149 3214 150
rect 3682 508 3688 511
rect 3682 504 3683 508
rect 3687 504 3688 508
rect 3682 502 3688 504
rect 3682 498 3683 502
rect 3687 498 3688 502
rect 3682 496 3688 498
rect 3682 492 3683 496
rect 3687 492 3688 496
rect 3682 490 3688 492
rect 3682 486 3683 490
rect 3687 486 3688 490
rect 3682 484 3688 486
rect 3682 480 3683 484
rect 3687 480 3688 484
rect 3682 478 3688 480
rect 3682 474 3683 478
rect 3687 474 3688 478
rect 3682 472 3688 474
rect 3682 468 3683 472
rect 3687 468 3688 472
rect 3682 466 3688 468
rect 3682 462 3683 466
rect 3687 462 3688 466
rect 3682 460 3688 462
rect 3682 456 3683 460
rect 3687 456 3688 460
rect 3682 454 3688 456
rect 3682 450 3683 454
rect 3687 450 3688 454
rect 3682 448 3688 450
rect 3682 444 3683 448
rect 3687 444 3688 448
rect 3682 442 3688 444
rect 3682 438 3683 442
rect 3687 438 3688 442
rect 3682 436 3688 438
rect 3682 432 3683 436
rect 3687 432 3688 436
rect 3682 430 3688 432
rect 3682 426 3683 430
rect 3687 426 3688 430
rect 3682 424 3688 426
rect 3682 420 3683 424
rect 3687 420 3688 424
rect 3682 418 3688 420
rect 3682 414 3683 418
rect 3687 414 3688 418
rect 3682 412 3688 414
rect 3682 408 3683 412
rect 3687 408 3688 412
rect 3682 406 3688 408
rect 3682 402 3683 406
rect 3687 402 3688 406
rect 3682 400 3688 402
rect 3682 396 3683 400
rect 3687 396 3688 400
rect 3682 394 3688 396
rect 3682 390 3683 394
rect 3687 390 3688 394
rect 3682 388 3688 390
rect 3682 384 3683 388
rect 3687 384 3688 388
rect 3682 382 3688 384
rect 3682 378 3683 382
rect 3687 378 3688 382
rect 3682 376 3688 378
rect 3682 372 3683 376
rect 3687 372 3688 376
rect 3682 370 3688 372
rect 3682 366 3683 370
rect 3687 366 3688 370
rect 3682 364 3688 366
rect 3682 360 3683 364
rect 3687 360 3688 364
rect 3682 358 3688 360
rect 3682 354 3683 358
rect 3687 354 3688 358
rect 3682 352 3688 354
rect 3682 348 3683 352
rect 3687 348 3688 352
rect 3682 346 3688 348
rect 3682 342 3683 346
rect 3687 342 3688 346
rect 3682 340 3688 342
rect 3682 336 3683 340
rect 3687 336 3688 340
rect 3682 334 3688 336
rect 3682 330 3683 334
rect 3687 330 3688 334
rect 3682 328 3688 330
rect 3682 324 3683 328
rect 3687 324 3688 328
rect 3682 322 3688 324
rect 3682 318 3683 322
rect 3687 318 3688 322
rect 3682 316 3688 318
rect 3682 312 3683 316
rect 3687 312 3688 316
rect 3682 310 3688 312
rect 3682 306 3683 310
rect 3687 306 3688 310
rect 3682 304 3688 306
rect 3682 300 3683 304
rect 3687 300 3688 304
rect 3682 298 3688 300
rect 3682 294 3683 298
rect 3687 294 3688 298
rect 3682 292 3688 294
rect 3682 288 3683 292
rect 3687 288 3688 292
rect 3682 286 3688 288
rect 3682 282 3683 286
rect 3687 282 3688 286
rect 3682 280 3688 282
rect 3682 276 3683 280
rect 3687 276 3688 280
rect 3682 274 3688 276
rect 3682 270 3683 274
rect 3687 270 3688 274
rect 3682 268 3688 270
rect 3682 264 3683 268
rect 3687 264 3688 268
rect 3682 262 3688 264
rect 3682 258 3683 262
rect 3687 258 3688 262
rect 3682 256 3688 258
rect 3682 252 3683 256
rect 3687 252 3688 256
rect 3682 250 3688 252
rect 3682 246 3683 250
rect 3687 246 3688 250
rect 3682 244 3688 246
rect 3682 240 3683 244
rect 3687 240 3688 244
rect 3682 238 3688 240
rect 3682 234 3683 238
rect 3687 234 3688 238
rect 3682 232 3688 234
rect 3682 228 3683 232
rect 3687 228 3688 232
rect 3682 226 3688 228
rect 3682 222 3683 226
rect 3687 222 3688 226
rect 3682 220 3688 222
rect 3682 216 3683 220
rect 3687 216 3688 220
rect 3682 214 3688 216
rect 3682 210 3683 214
rect 3687 210 3688 214
rect 3682 208 3688 210
rect 3682 204 3683 208
rect 3687 204 3688 208
rect 3682 202 3688 204
rect 3682 198 3683 202
rect 3687 198 3688 202
rect 3682 196 3688 198
rect 3682 192 3683 196
rect 3687 192 3688 196
rect 3682 190 3688 192
rect 3682 186 3683 190
rect 3687 186 3688 190
rect 3682 184 3688 186
rect 3682 180 3683 184
rect 3687 180 3688 184
rect 3682 178 3688 180
rect 3682 174 3683 178
rect 3687 174 3688 178
rect 3682 172 3688 174
rect 3682 168 3683 172
rect 3687 168 3688 172
rect 3682 166 3688 168
rect 3682 162 3683 166
rect 3687 162 3688 166
rect 3682 160 3688 162
rect 3682 156 3683 160
rect 3687 156 3688 160
rect 3682 154 3688 156
rect 3682 150 3683 154
rect 3687 150 3688 154
rect 3682 149 3688 150
rect 4156 508 4162 511
rect 4156 504 4157 508
rect 4161 504 4162 508
rect 4156 502 4162 504
rect 4156 498 4157 502
rect 4161 498 4162 502
rect 4156 496 4162 498
rect 4156 492 4157 496
rect 4161 492 4162 496
rect 4156 490 4162 492
rect 4156 486 4157 490
rect 4161 486 4162 490
rect 4156 484 4162 486
rect 4156 480 4157 484
rect 4161 480 4162 484
rect 4156 478 4162 480
rect 4156 474 4157 478
rect 4161 474 4162 478
rect 4156 472 4162 474
rect 4156 468 4157 472
rect 4161 468 4162 472
rect 4156 466 4162 468
rect 4156 462 4157 466
rect 4161 462 4162 466
rect 4156 460 4162 462
rect 4156 456 4157 460
rect 4161 456 4162 460
rect 4156 454 4162 456
rect 4156 450 4157 454
rect 4161 450 4162 454
rect 4156 448 4162 450
rect 4156 444 4157 448
rect 4161 444 4162 448
rect 4156 442 4162 444
rect 4156 438 4157 442
rect 4161 438 4162 442
rect 4156 436 4162 438
rect 4156 432 4157 436
rect 4161 432 4162 436
rect 4156 430 4162 432
rect 4156 426 4157 430
rect 4161 426 4162 430
rect 4156 424 4162 426
rect 4156 420 4157 424
rect 4161 420 4162 424
rect 4156 418 4162 420
rect 4156 414 4157 418
rect 4161 414 4162 418
rect 4156 412 4162 414
rect 4156 408 4157 412
rect 4161 408 4162 412
rect 4156 406 4162 408
rect 4156 402 4157 406
rect 4161 402 4162 406
rect 4156 400 4162 402
rect 4156 396 4157 400
rect 4161 396 4162 400
rect 4156 394 4162 396
rect 4156 390 4157 394
rect 4161 390 4162 394
rect 4156 388 4162 390
rect 4156 384 4157 388
rect 4161 384 4162 388
rect 4156 382 4162 384
rect 4156 378 4157 382
rect 4161 378 4162 382
rect 4156 376 4162 378
rect 4156 372 4157 376
rect 4161 372 4162 376
rect 4156 370 4162 372
rect 4156 366 4157 370
rect 4161 366 4162 370
rect 4156 364 4162 366
rect 4156 360 4157 364
rect 4161 360 4162 364
rect 4156 358 4162 360
rect 4156 354 4157 358
rect 4161 354 4162 358
rect 4156 352 4162 354
rect 4156 348 4157 352
rect 4161 348 4162 352
rect 4156 346 4162 348
rect 4156 342 4157 346
rect 4161 342 4162 346
rect 4156 340 4162 342
rect 4156 336 4157 340
rect 4161 336 4162 340
rect 4156 334 4162 336
rect 4156 330 4157 334
rect 4161 330 4162 334
rect 4156 328 4162 330
rect 4156 324 4157 328
rect 4161 324 4162 328
rect 4156 322 4162 324
rect 4156 318 4157 322
rect 4161 318 4162 322
rect 4156 316 4162 318
rect 4156 312 4157 316
rect 4161 312 4162 316
rect 4156 310 4162 312
rect 4156 306 4157 310
rect 4161 306 4162 310
rect 4156 304 4162 306
rect 4156 300 4157 304
rect 4161 300 4162 304
rect 4156 298 4162 300
rect 4156 294 4157 298
rect 4161 294 4162 298
rect 4156 292 4162 294
rect 4156 288 4157 292
rect 4161 288 4162 292
rect 4156 286 4162 288
rect 4156 282 4157 286
rect 4161 282 4162 286
rect 4156 280 4162 282
rect 4156 276 4157 280
rect 4161 276 4162 280
rect 4156 274 4162 276
rect 4156 270 4157 274
rect 4161 270 4162 274
rect 4156 268 4162 270
rect 4156 264 4157 268
rect 4161 264 4162 268
rect 4156 262 4162 264
rect 4156 258 4157 262
rect 4161 258 4162 262
rect 4156 256 4162 258
rect 4156 252 4157 256
rect 4161 252 4162 256
rect 4156 250 4162 252
rect 4156 246 4157 250
rect 4161 246 4162 250
rect 4156 244 4162 246
rect 4156 240 4157 244
rect 4161 240 4162 244
rect 4156 238 4162 240
rect 4156 234 4157 238
rect 4161 234 4162 238
rect 4156 232 4162 234
rect 4156 228 4157 232
rect 4161 228 4162 232
rect 4156 226 4162 228
rect 4156 222 4157 226
rect 4161 222 4162 226
rect 4156 220 4162 222
rect 4156 216 4157 220
rect 4161 216 4162 220
rect 4156 214 4162 216
rect 4156 210 4157 214
rect 4161 210 4162 214
rect 4156 208 4162 210
rect 4156 204 4157 208
rect 4161 204 4162 208
rect 4156 202 4162 204
rect 4156 198 4157 202
rect 4161 198 4162 202
rect 4156 196 4162 198
rect 4156 192 4157 196
rect 4161 192 4162 196
rect 4156 190 4162 192
rect 4156 186 4157 190
rect 4161 186 4162 190
rect 4156 184 4162 186
rect 4156 180 4157 184
rect 4161 180 4162 184
rect 4156 178 4162 180
rect 4156 174 4157 178
rect 4161 174 4162 178
rect 4156 172 4162 174
rect 4156 168 4157 172
rect 4161 168 4162 172
rect 4156 166 4162 168
rect 4156 162 4157 166
rect 4161 162 4162 166
rect 4156 160 4162 162
rect 4156 156 4157 160
rect 4161 156 4162 160
rect 4156 154 4162 156
rect 4156 150 4157 154
rect 4161 150 4162 154
rect 4156 149 4162 150
rect 4630 508 4636 511
rect 4630 504 4631 508
rect 4635 504 4636 508
rect 4630 502 4636 504
rect 4630 498 4631 502
rect 4635 498 4636 502
rect 4630 496 4636 498
rect 4630 492 4631 496
rect 4635 492 4636 496
rect 4630 490 4636 492
rect 4630 486 4631 490
rect 4635 486 4636 490
rect 4630 484 4636 486
rect 4630 480 4631 484
rect 4635 480 4636 484
rect 4630 478 4636 480
rect 4630 474 4631 478
rect 4635 474 4636 478
rect 4630 472 4636 474
rect 4630 468 4631 472
rect 4635 468 4636 472
rect 4630 466 4636 468
rect 4630 462 4631 466
rect 4635 462 4636 466
rect 4630 460 4636 462
rect 4630 456 4631 460
rect 4635 456 4636 460
rect 4630 454 4636 456
rect 4630 450 4631 454
rect 4635 450 4636 454
rect 4630 448 4636 450
rect 4630 444 4631 448
rect 4635 444 4636 448
rect 4630 442 4636 444
rect 4630 438 4631 442
rect 4635 438 4636 442
rect 4630 436 4636 438
rect 4630 432 4631 436
rect 4635 432 4636 436
rect 4630 430 4636 432
rect 4630 426 4631 430
rect 4635 426 4636 430
rect 4630 424 4636 426
rect 4630 420 4631 424
rect 4635 420 4636 424
rect 4630 418 4636 420
rect 4630 414 4631 418
rect 4635 414 4636 418
rect 4630 412 4636 414
rect 4630 408 4631 412
rect 4635 408 4636 412
rect 4630 406 4636 408
rect 4630 402 4631 406
rect 4635 402 4636 406
rect 4630 400 4636 402
rect 4630 396 4631 400
rect 4635 396 4636 400
rect 4630 394 4636 396
rect 4630 390 4631 394
rect 4635 390 4636 394
rect 4630 388 4636 390
rect 4630 384 4631 388
rect 4635 384 4636 388
rect 4630 382 4636 384
rect 4630 378 4631 382
rect 4635 378 4636 382
rect 4630 376 4636 378
rect 4630 372 4631 376
rect 4635 372 4636 376
rect 4630 370 4636 372
rect 4630 366 4631 370
rect 4635 366 4636 370
rect 4630 364 4636 366
rect 4630 360 4631 364
rect 4635 360 4636 364
rect 4630 358 4636 360
rect 4630 354 4631 358
rect 4635 354 4636 358
rect 4630 352 4636 354
rect 4630 348 4631 352
rect 4635 348 4636 352
rect 4630 346 4636 348
rect 4630 342 4631 346
rect 4635 342 4636 346
rect 4630 340 4636 342
rect 4630 336 4631 340
rect 4635 336 4636 340
rect 4630 334 4636 336
rect 4630 330 4631 334
rect 4635 330 4636 334
rect 4630 328 4636 330
rect 4630 324 4631 328
rect 4635 324 4636 328
rect 4630 322 4636 324
rect 4630 318 4631 322
rect 4635 318 4636 322
rect 4630 316 4636 318
rect 4630 312 4631 316
rect 4635 312 4636 316
rect 4630 310 4636 312
rect 4630 306 4631 310
rect 4635 306 4636 310
rect 4630 304 4636 306
rect 4630 300 4631 304
rect 4635 300 4636 304
rect 4630 298 4636 300
rect 4630 294 4631 298
rect 4635 294 4636 298
rect 4630 292 4636 294
rect 4630 288 4631 292
rect 4635 288 4636 292
rect 4630 286 4636 288
rect 4630 282 4631 286
rect 4635 282 4636 286
rect 4630 280 4636 282
rect 4630 276 4631 280
rect 4635 276 4636 280
rect 4630 274 4636 276
rect 4630 270 4631 274
rect 4635 270 4636 274
rect 4630 268 4636 270
rect 4630 264 4631 268
rect 4635 264 4636 268
rect 4630 262 4636 264
rect 4630 258 4631 262
rect 4635 258 4636 262
rect 4630 256 4636 258
rect 4630 252 4631 256
rect 4635 252 4636 256
rect 4630 250 4636 252
rect 4630 246 4631 250
rect 4635 246 4636 250
rect 4630 244 4636 246
rect 4630 240 4631 244
rect 4635 240 4636 244
rect 4630 238 4636 240
rect 4630 234 4631 238
rect 4635 234 4636 238
rect 4630 232 4636 234
rect 4630 228 4631 232
rect 4635 228 4636 232
rect 4630 226 4636 228
rect 4630 222 4631 226
rect 4635 222 4636 226
rect 4630 220 4636 222
rect 4630 216 4631 220
rect 4635 216 4636 220
rect 4630 214 4636 216
rect 4630 210 4631 214
rect 4635 210 4636 214
rect 4630 208 4636 210
rect 4630 204 4631 208
rect 4635 204 4636 208
rect 4630 202 4636 204
rect 4630 198 4631 202
rect 4635 199 4636 202
rect 4635 198 4800 199
rect 4630 196 4800 198
rect 4630 192 4631 196
rect 4635 193 4800 196
rect 4635 192 4636 193
rect 4630 190 4636 192
rect 4630 186 4631 190
rect 4635 186 4636 190
rect 4630 184 4636 186
rect 4630 180 4631 184
rect 4635 180 4636 184
rect 4630 178 4636 180
rect 4630 174 4631 178
rect 4635 174 4636 178
rect 4630 172 4636 174
rect 4630 168 4631 172
rect 4635 168 4636 172
rect 4630 166 4636 168
rect 4630 162 4631 166
rect 4635 162 4636 166
rect 4630 160 4636 162
rect 4630 156 4631 160
rect 4635 156 4636 160
rect 4630 154 4636 156
rect 4686 186 4692 193
rect 4686 182 4687 186
rect 4691 182 4692 186
rect 4686 180 4692 182
rect 4686 176 4687 180
rect 4691 176 4692 180
rect 4686 174 4692 176
rect 4686 170 4687 174
rect 4691 170 4692 174
rect 4686 168 4692 170
rect 4686 164 4687 168
rect 4691 164 4692 168
rect 4686 162 4692 164
rect 4686 158 4687 162
rect 4691 158 4692 162
rect 4686 156 4692 158
rect 4630 150 4631 154
rect 4635 150 4636 154
rect 4630 149 4636 150
rect 4686 152 4687 156
rect 4691 152 4692 156
rect 4742 186 4748 193
rect 4742 182 4743 186
rect 4747 182 4748 186
rect 4742 180 4748 182
rect 4742 176 4743 180
rect 4747 176 4748 180
rect 4742 174 4748 176
rect 4742 170 4743 174
rect 4747 170 4748 174
rect 4742 168 4748 170
rect 4742 164 4743 168
rect 4747 164 4748 168
rect 4742 162 4748 164
rect 4742 158 4743 162
rect 4747 158 4748 162
rect 4742 156 4748 158
rect 4686 149 4692 152
rect 4742 152 4743 156
rect 4747 152 4748 156
rect 4768 186 4774 193
rect 4768 182 4769 186
rect 4773 182 4774 186
rect 4768 180 4774 182
rect 4768 176 4769 180
rect 4773 176 4774 180
rect 4768 174 4774 176
rect 4768 170 4769 174
rect 4773 170 4774 174
rect 4768 168 4774 170
rect 4768 164 4769 168
rect 4773 164 4774 168
rect 4768 162 4774 164
rect 4768 158 4769 162
rect 4773 158 4774 162
rect 4768 156 4774 158
rect 4742 149 4748 152
rect 4768 152 4769 156
rect 4773 152 4774 156
rect 4794 186 4800 193
rect 4794 182 4795 186
rect 4799 182 4800 186
rect 4794 180 4800 182
rect 4794 176 4795 180
rect 4799 176 4800 180
rect 4794 174 4800 176
rect 4794 170 4795 174
rect 4799 170 4800 174
rect 4794 168 4800 170
rect 4794 164 4795 168
rect 4799 164 4800 168
rect 4794 162 4800 164
rect 4794 158 4795 162
rect 4799 158 4800 162
rect 4794 156 4800 158
rect 4768 149 4774 152
rect 4794 152 4795 156
rect 4799 152 4800 156
rect 4794 149 4800 152
rect 2 148 4998 149
rect 2 144 5 148
rect 9 144 11 148
rect 15 144 17 148
rect 21 144 23 148
rect 27 144 29 148
rect 33 144 35 148
rect 39 144 41 148
rect 45 144 47 148
rect 51 144 53 148
rect 57 144 59 148
rect 63 144 65 148
rect 69 144 71 148
rect 75 144 77 148
rect 81 144 83 148
rect 87 144 89 148
rect 93 144 95 148
rect 99 144 101 148
rect 105 144 107 148
rect 111 144 113 148
rect 117 144 119 148
rect 123 144 125 148
rect 129 144 131 148
rect 135 144 137 148
rect 141 144 143 148
rect 147 144 149 148
rect 153 144 155 148
rect 159 144 161 148
rect 165 144 167 148
rect 171 144 173 148
rect 177 144 179 148
rect 183 144 185 148
rect 189 144 191 148
rect 195 144 197 148
rect 201 144 203 148
rect 207 144 209 148
rect 213 144 215 148
rect 219 144 221 148
rect 225 144 227 148
rect 231 144 233 148
rect 237 144 239 148
rect 243 144 245 148
rect 249 144 251 148
rect 255 144 257 148
rect 261 144 263 148
rect 267 144 269 148
rect 273 144 275 148
rect 279 144 281 148
rect 285 144 287 148
rect 291 144 293 148
rect 297 144 299 148
rect 303 144 305 148
rect 309 144 311 148
rect 315 144 317 148
rect 321 144 323 148
rect 327 144 329 148
rect 333 144 335 148
rect 339 144 341 148
rect 345 144 347 148
rect 351 144 353 148
rect 357 144 359 148
rect 363 144 365 148
rect 369 144 371 148
rect 375 144 377 148
rect 381 144 383 148
rect 387 144 389 148
rect 393 144 395 148
rect 399 144 401 148
rect 405 144 407 148
rect 411 144 413 148
rect 417 144 419 148
rect 423 144 425 148
rect 429 144 431 148
rect 435 144 437 148
rect 441 144 443 148
rect 447 144 449 148
rect 453 144 455 148
rect 459 144 461 148
rect 465 144 467 148
rect 471 144 473 148
rect 477 144 479 148
rect 483 144 485 148
rect 489 144 491 148
rect 495 144 497 148
rect 501 144 503 148
rect 507 144 509 148
rect 513 144 515 148
rect 519 144 521 148
rect 525 144 527 148
rect 531 144 533 148
rect 537 144 539 148
rect 543 144 545 148
rect 549 144 551 148
rect 555 144 557 148
rect 561 144 563 148
rect 567 144 569 148
rect 573 144 575 148
rect 579 144 581 148
rect 585 144 587 148
rect 591 144 617 148
rect 621 144 623 148
rect 627 144 629 148
rect 633 144 635 148
rect 639 144 641 148
rect 645 144 647 148
rect 651 144 653 148
rect 657 144 659 148
rect 663 144 665 148
rect 669 144 671 148
rect 675 144 677 148
rect 681 144 683 148
rect 687 144 689 148
rect 693 144 695 148
rect 699 144 701 148
rect 705 144 707 148
rect 711 144 713 148
rect 717 144 719 148
rect 723 144 725 148
rect 729 144 731 148
rect 735 144 737 148
rect 741 144 743 148
rect 747 144 749 148
rect 753 144 755 148
rect 759 144 761 148
rect 765 144 767 148
rect 771 144 773 148
rect 777 144 779 148
rect 783 144 785 148
rect 789 144 791 148
rect 795 144 797 148
rect 801 144 803 148
rect 807 144 809 148
rect 813 144 815 148
rect 819 144 821 148
rect 825 144 827 148
rect 831 144 833 148
rect 837 144 839 148
rect 843 144 845 148
rect 849 144 851 148
rect 855 144 857 148
rect 861 144 863 148
rect 867 144 869 148
rect 873 144 875 148
rect 879 144 881 148
rect 885 144 887 148
rect 891 144 893 148
rect 897 144 899 148
rect 903 144 905 148
rect 909 144 911 148
rect 915 144 917 148
rect 921 144 923 148
rect 927 144 929 148
rect 933 144 935 148
rect 939 144 941 148
rect 945 144 947 148
rect 951 144 953 148
rect 957 144 959 148
rect 963 144 965 148
rect 969 144 971 148
rect 975 144 977 148
rect 981 144 983 148
rect 987 144 989 148
rect 993 144 995 148
rect 999 144 1001 148
rect 1005 144 1007 148
rect 1011 144 1013 148
rect 1017 144 1019 148
rect 1023 144 1025 148
rect 1029 144 1031 148
rect 1035 144 1037 148
rect 1041 144 1043 148
rect 1047 144 1049 148
rect 1053 144 1055 148
rect 1059 144 1061 148
rect 1065 144 1091 148
rect 1095 144 1097 148
rect 1101 144 1103 148
rect 1107 144 1109 148
rect 1113 144 1115 148
rect 1119 144 1121 148
rect 1125 144 1127 148
rect 1131 144 1133 148
rect 1137 144 1139 148
rect 1143 144 1145 148
rect 1149 144 1151 148
rect 1155 144 1157 148
rect 1161 144 1163 148
rect 1167 144 1169 148
rect 1173 144 1175 148
rect 1179 144 1181 148
rect 1185 144 1187 148
rect 1191 144 1193 148
rect 1197 144 1199 148
rect 1203 144 1205 148
rect 1209 144 1211 148
rect 1215 144 1217 148
rect 1221 144 1223 148
rect 1227 144 1229 148
rect 1233 144 1235 148
rect 1239 144 1241 148
rect 1245 144 1247 148
rect 1251 144 1253 148
rect 1257 144 1259 148
rect 1263 144 1265 148
rect 1269 144 1271 148
rect 1275 144 1277 148
rect 1281 144 1283 148
rect 1287 144 1289 148
rect 1293 144 1295 148
rect 1299 144 1301 148
rect 1305 144 1307 148
rect 1311 144 1313 148
rect 1317 144 1319 148
rect 1323 144 1325 148
rect 1329 144 1331 148
rect 1335 144 1337 148
rect 1341 144 1343 148
rect 1347 144 1349 148
rect 1353 144 1355 148
rect 1359 144 1361 148
rect 1365 144 1367 148
rect 1371 144 1373 148
rect 1377 144 1379 148
rect 1383 144 1385 148
rect 1389 144 1391 148
rect 1395 144 1397 148
rect 1401 144 1403 148
rect 1407 144 1409 148
rect 1413 144 1415 148
rect 1419 144 1421 148
rect 1425 144 1427 148
rect 1431 144 1433 148
rect 1437 144 1439 148
rect 1443 144 1445 148
rect 1449 144 1451 148
rect 1455 144 1457 148
rect 1461 144 1463 148
rect 1467 144 1469 148
rect 1473 144 1475 148
rect 1479 144 1481 148
rect 1485 144 1487 148
rect 1491 144 1493 148
rect 1497 144 1499 148
rect 1503 144 1505 148
rect 1509 144 1511 148
rect 1515 144 1517 148
rect 1521 144 1523 148
rect 1527 144 1529 148
rect 1533 144 1535 148
rect 1539 144 1565 148
rect 1569 144 1571 148
rect 1575 144 1577 148
rect 1581 144 1583 148
rect 1587 144 1589 148
rect 1593 144 1595 148
rect 1599 144 1601 148
rect 1605 144 1607 148
rect 1611 144 1613 148
rect 1617 144 1619 148
rect 1623 144 1625 148
rect 1629 144 1631 148
rect 1635 144 1637 148
rect 1641 144 1643 148
rect 1647 144 1649 148
rect 1653 144 1655 148
rect 1659 144 1661 148
rect 1665 144 1667 148
rect 1671 144 1673 148
rect 1677 144 1679 148
rect 1683 144 1685 148
rect 1689 144 1691 148
rect 1695 144 1697 148
rect 1701 144 1703 148
rect 1707 144 1709 148
rect 1713 144 1715 148
rect 1719 144 1721 148
rect 1725 144 1727 148
rect 1731 144 1733 148
rect 1737 144 1739 148
rect 1743 144 1745 148
rect 1749 144 1751 148
rect 1755 144 1757 148
rect 1761 144 1763 148
rect 1767 144 1769 148
rect 1773 144 1775 148
rect 1779 144 1781 148
rect 1785 144 1787 148
rect 1791 144 1793 148
rect 1797 144 1799 148
rect 1803 144 1805 148
rect 1809 144 1811 148
rect 1815 144 1817 148
rect 1821 144 1823 148
rect 1827 144 1829 148
rect 1833 144 1835 148
rect 1839 144 1841 148
rect 1845 144 1847 148
rect 1851 144 1853 148
rect 1857 144 1859 148
rect 1863 144 1865 148
rect 1869 144 1871 148
rect 1875 144 1877 148
rect 1881 144 1883 148
rect 1887 144 1889 148
rect 1893 144 1895 148
rect 1899 144 1901 148
rect 1905 144 1907 148
rect 1911 144 1913 148
rect 1917 144 1919 148
rect 1923 144 1925 148
rect 1929 144 1931 148
rect 1935 144 1937 148
rect 1941 144 1943 148
rect 1947 144 1949 148
rect 1953 144 1955 148
rect 1959 144 1961 148
rect 1965 144 1967 148
rect 1971 144 1973 148
rect 1977 144 1979 148
rect 1983 144 1985 148
rect 1989 144 1991 148
rect 1995 144 1997 148
rect 2001 144 2003 148
rect 2007 144 2009 148
rect 2013 144 2039 148
rect 2043 144 2045 148
rect 2049 144 2051 148
rect 2055 144 2057 148
rect 2061 144 2063 148
rect 2067 144 2069 148
rect 2073 144 2075 148
rect 2079 144 2081 148
rect 2085 144 2087 148
rect 2091 144 2093 148
rect 2097 144 2099 148
rect 2103 144 2105 148
rect 2109 144 2111 148
rect 2115 144 2117 148
rect 2121 144 2123 148
rect 2127 144 2129 148
rect 2133 144 2135 148
rect 2139 144 2141 148
rect 2145 144 2147 148
rect 2151 144 2153 148
rect 2157 144 2159 148
rect 2163 144 2165 148
rect 2169 144 2171 148
rect 2175 144 2177 148
rect 2181 144 2183 148
rect 2187 144 2189 148
rect 2193 144 2195 148
rect 2199 144 2201 148
rect 2205 144 2207 148
rect 2211 144 2213 148
rect 2217 144 2219 148
rect 2223 144 2225 148
rect 2229 144 2231 148
rect 2235 144 2237 148
rect 2241 144 2243 148
rect 2247 144 2249 148
rect 2253 144 2255 148
rect 2259 144 2261 148
rect 2265 144 2267 148
rect 2271 144 2273 148
rect 2277 144 2279 148
rect 2283 144 2285 148
rect 2289 144 2291 148
rect 2295 144 2297 148
rect 2301 144 2303 148
rect 2307 144 2309 148
rect 2313 144 2315 148
rect 2319 144 2321 148
rect 2325 144 2327 148
rect 2331 144 2333 148
rect 2337 144 2339 148
rect 2343 144 2345 148
rect 2349 144 2351 148
rect 2355 144 2357 148
rect 2361 144 2363 148
rect 2367 144 2369 148
rect 2373 144 2375 148
rect 2379 144 2381 148
rect 2385 144 2387 148
rect 2391 144 2393 148
rect 2397 144 2399 148
rect 2403 144 2405 148
rect 2409 144 2411 148
rect 2415 144 2417 148
rect 2421 144 2423 148
rect 2427 144 2429 148
rect 2433 144 2435 148
rect 2439 144 2441 148
rect 2445 144 2447 148
rect 2451 144 2453 148
rect 2457 144 2459 148
rect 2463 144 2465 148
rect 2469 144 2471 148
rect 2475 144 2477 148
rect 2481 144 2483 148
rect 2487 144 2513 148
rect 2517 144 2519 148
rect 2523 144 2525 148
rect 2529 144 2531 148
rect 2535 144 2537 148
rect 2541 144 2543 148
rect 2547 144 2549 148
rect 2553 144 2555 148
rect 2559 144 2561 148
rect 2565 144 2567 148
rect 2571 144 2573 148
rect 2577 144 2579 148
rect 2583 144 2585 148
rect 2589 144 2591 148
rect 2595 144 2597 148
rect 2601 144 2603 148
rect 2607 144 2609 148
rect 2613 144 2615 148
rect 2619 144 2621 148
rect 2625 144 2627 148
rect 2631 144 2633 148
rect 2637 144 2639 148
rect 2643 144 2645 148
rect 2649 144 2651 148
rect 2655 144 2657 148
rect 2661 144 2663 148
rect 2667 144 2669 148
rect 2673 144 2675 148
rect 2679 144 2681 148
rect 2685 144 2687 148
rect 2691 144 2693 148
rect 2697 144 2699 148
rect 2703 144 2705 148
rect 2709 144 2711 148
rect 2715 144 2717 148
rect 2721 144 2723 148
rect 2727 144 2729 148
rect 2733 144 2735 148
rect 2739 144 2741 148
rect 2745 144 2747 148
rect 2751 144 2753 148
rect 2757 144 2759 148
rect 2763 144 2765 148
rect 2769 144 2771 148
rect 2775 144 2777 148
rect 2781 144 2783 148
rect 2787 144 2789 148
rect 2793 144 2795 148
rect 2799 144 2801 148
rect 2805 144 2807 148
rect 2811 144 2813 148
rect 2817 144 2819 148
rect 2823 144 2825 148
rect 2829 144 2831 148
rect 2835 144 2837 148
rect 2841 144 2843 148
rect 2847 144 2849 148
rect 2853 144 2855 148
rect 2859 144 2861 148
rect 2865 144 2867 148
rect 2871 144 2873 148
rect 2877 144 2879 148
rect 2883 144 2885 148
rect 2889 144 2891 148
rect 2895 144 2897 148
rect 2901 144 2903 148
rect 2907 144 2909 148
rect 2913 144 2915 148
rect 2919 144 2921 148
rect 2925 144 2927 148
rect 2931 144 2933 148
rect 2937 144 2939 148
rect 2943 144 2945 148
rect 2949 144 2951 148
rect 2955 144 2957 148
rect 2961 144 2987 148
rect 2991 144 2993 148
rect 2997 144 2999 148
rect 3003 144 3005 148
rect 3009 144 3011 148
rect 3015 144 3017 148
rect 3021 144 3023 148
rect 3027 144 3029 148
rect 3033 144 3035 148
rect 3039 144 3041 148
rect 3045 144 3047 148
rect 3051 144 3053 148
rect 3057 144 3059 148
rect 3063 144 3065 148
rect 3069 144 3071 148
rect 3075 144 3077 148
rect 3081 144 3083 148
rect 3087 144 3089 148
rect 3093 144 3095 148
rect 3099 144 3101 148
rect 3105 144 3107 148
rect 3111 144 3113 148
rect 3117 144 3119 148
rect 3123 144 3125 148
rect 3129 144 3131 148
rect 3135 144 3137 148
rect 3141 144 3143 148
rect 3147 144 3149 148
rect 3153 144 3155 148
rect 3159 144 3161 148
rect 3165 144 3167 148
rect 3171 144 3173 148
rect 3177 144 3179 148
rect 3183 144 3185 148
rect 3189 144 3191 148
rect 3195 144 3197 148
rect 3201 144 3203 148
rect 3207 144 3209 148
rect 3213 144 3215 148
rect 3219 144 3221 148
rect 3225 144 3227 148
rect 3231 144 3233 148
rect 3237 144 3239 148
rect 3243 144 3245 148
rect 3249 144 3251 148
rect 3255 144 3257 148
rect 3261 144 3263 148
rect 3267 144 3269 148
rect 3273 144 3275 148
rect 3279 144 3281 148
rect 3285 144 3287 148
rect 3291 144 3293 148
rect 3297 144 3299 148
rect 3303 144 3305 148
rect 3309 144 3311 148
rect 3315 144 3317 148
rect 3321 144 3323 148
rect 3327 144 3329 148
rect 3333 144 3335 148
rect 3339 144 3341 148
rect 3345 144 3347 148
rect 3351 144 3353 148
rect 3357 144 3359 148
rect 3363 144 3365 148
rect 3369 144 3371 148
rect 3375 144 3377 148
rect 3381 144 3383 148
rect 3387 144 3389 148
rect 3393 144 3395 148
rect 3399 144 3401 148
rect 3405 144 3407 148
rect 3411 144 3413 148
rect 3417 144 3419 148
rect 3423 144 3425 148
rect 3429 144 3431 148
rect 3435 144 3461 148
rect 3465 144 3467 148
rect 3471 144 3473 148
rect 3477 144 3479 148
rect 3483 144 3485 148
rect 3489 144 3491 148
rect 3495 144 3497 148
rect 3501 144 3503 148
rect 3507 144 3509 148
rect 3513 144 3515 148
rect 3519 144 3521 148
rect 3525 144 3527 148
rect 3531 144 3533 148
rect 3537 144 3539 148
rect 3543 144 3545 148
rect 3549 144 3551 148
rect 3555 144 3557 148
rect 3561 144 3563 148
rect 3567 144 3569 148
rect 3573 144 3575 148
rect 3579 144 3581 148
rect 3585 144 3587 148
rect 3591 144 3593 148
rect 3597 144 3599 148
rect 3603 144 3605 148
rect 3609 144 3611 148
rect 3615 144 3617 148
rect 3621 144 3623 148
rect 3627 144 3629 148
rect 3633 144 3635 148
rect 3639 144 3641 148
rect 3645 144 3647 148
rect 3651 144 3653 148
rect 3657 144 3659 148
rect 3663 144 3665 148
rect 3669 144 3671 148
rect 3675 144 3677 148
rect 3681 144 3683 148
rect 3687 144 3689 148
rect 3693 144 3695 148
rect 3699 144 3701 148
rect 3705 144 3707 148
rect 3711 144 3713 148
rect 3717 144 3719 148
rect 3723 144 3725 148
rect 3729 144 3731 148
rect 3735 144 3737 148
rect 3741 144 3743 148
rect 3747 144 3749 148
rect 3753 144 3755 148
rect 3759 144 3761 148
rect 3765 144 3767 148
rect 3771 144 3773 148
rect 3777 144 3779 148
rect 3783 144 3785 148
rect 3789 144 3791 148
rect 3795 144 3797 148
rect 3801 144 3803 148
rect 3807 144 3809 148
rect 3813 144 3815 148
rect 3819 144 3821 148
rect 3825 144 3827 148
rect 3831 144 3833 148
rect 3837 144 3839 148
rect 3843 144 3845 148
rect 3849 144 3851 148
rect 3855 144 3857 148
rect 3861 144 3863 148
rect 3867 144 3869 148
rect 3873 144 3875 148
rect 3879 144 3881 148
rect 3885 144 3887 148
rect 3891 144 3893 148
rect 3897 144 3899 148
rect 3903 144 3905 148
rect 3909 144 3935 148
rect 3939 144 3941 148
rect 3945 144 3947 148
rect 3951 144 3953 148
rect 3957 144 3959 148
rect 3963 144 3965 148
rect 3969 144 3971 148
rect 3975 144 3977 148
rect 3981 144 3983 148
rect 3987 144 3989 148
rect 3993 144 3995 148
rect 3999 144 4001 148
rect 4005 144 4007 148
rect 4011 144 4013 148
rect 4017 144 4019 148
rect 4023 144 4025 148
rect 4029 144 4031 148
rect 4035 144 4037 148
rect 4041 144 4043 148
rect 4047 144 4049 148
rect 4053 144 4055 148
rect 4059 144 4061 148
rect 4065 144 4067 148
rect 4071 144 4073 148
rect 4077 144 4079 148
rect 4083 144 4085 148
rect 4089 144 4091 148
rect 4095 144 4097 148
rect 4101 144 4103 148
rect 4107 144 4109 148
rect 4113 144 4115 148
rect 4119 144 4121 148
rect 4125 144 4127 148
rect 4131 144 4133 148
rect 4137 144 4139 148
rect 4143 144 4145 148
rect 4149 144 4151 148
rect 4155 144 4157 148
rect 4161 144 4163 148
rect 4167 144 4169 148
rect 4173 144 4175 148
rect 4179 144 4181 148
rect 4185 144 4187 148
rect 4191 144 4193 148
rect 4197 144 4199 148
rect 4203 144 4205 148
rect 4209 144 4211 148
rect 4215 144 4217 148
rect 4221 144 4223 148
rect 4227 144 4229 148
rect 4233 144 4235 148
rect 4239 144 4241 148
rect 4245 144 4247 148
rect 4251 144 4253 148
rect 4257 144 4259 148
rect 4263 144 4265 148
rect 4269 144 4271 148
rect 4275 144 4277 148
rect 4281 144 4283 148
rect 4287 144 4289 148
rect 4293 144 4295 148
rect 4299 144 4301 148
rect 4305 144 4307 148
rect 4311 144 4313 148
rect 4317 144 4319 148
rect 4323 144 4325 148
rect 4329 144 4331 148
rect 4335 144 4337 148
rect 4341 144 4343 148
rect 4347 144 4349 148
rect 4353 144 4355 148
rect 4359 144 4361 148
rect 4365 144 4367 148
rect 4371 144 4373 148
rect 4377 144 4379 148
rect 4383 144 4409 148
rect 4413 144 4415 148
rect 4419 144 4421 148
rect 4425 144 4427 148
rect 4431 144 4433 148
rect 4437 144 4439 148
rect 4443 144 4445 148
rect 4449 144 4451 148
rect 4455 144 4457 148
rect 4461 144 4463 148
rect 4467 144 4469 148
rect 4473 144 4475 148
rect 4479 144 4481 148
rect 4485 144 4487 148
rect 4491 144 4493 148
rect 4497 144 4499 148
rect 4503 144 4505 148
rect 4509 144 4511 148
rect 4515 144 4517 148
rect 4521 144 4523 148
rect 4527 144 4529 148
rect 4533 144 4535 148
rect 4539 144 4541 148
rect 4545 144 4547 148
rect 4551 144 4553 148
rect 4557 144 4559 148
rect 4563 144 4565 148
rect 4569 144 4571 148
rect 4575 144 4577 148
rect 4581 144 4583 148
rect 4587 144 4589 148
rect 4593 144 4595 148
rect 4599 144 4601 148
rect 4605 144 4607 148
rect 4611 144 4613 148
rect 4617 144 4619 148
rect 4623 144 4625 148
rect 4629 144 4631 148
rect 4635 144 4637 148
rect 4641 144 4643 148
rect 4647 144 4649 148
rect 4653 144 4655 148
rect 4659 144 4661 148
rect 4665 144 4667 148
rect 4671 144 4673 148
rect 4677 144 4679 148
rect 4683 144 4685 148
rect 4689 144 4691 148
rect 4695 144 4697 148
rect 4701 144 4703 148
rect 4707 144 4709 148
rect 4713 144 4715 148
rect 4719 144 4721 148
rect 4725 144 4727 148
rect 4731 144 4733 148
rect 4737 144 4739 148
rect 4743 144 4745 148
rect 4749 144 4751 148
rect 4755 144 4757 148
rect 4761 144 4763 148
rect 4767 144 4769 148
rect 4773 144 4775 148
rect 4779 144 4781 148
rect 4785 144 4787 148
rect 4791 144 4793 148
rect 4797 144 4799 148
rect 4803 144 4805 148
rect 4809 144 4811 148
rect 4815 144 4817 148
rect 4821 144 4823 148
rect 4827 144 4829 148
rect 4833 144 4835 148
rect 4839 144 4841 148
rect 4845 144 4847 148
rect 4851 144 4853 148
rect 4857 144 4859 148
rect 4863 144 4865 148
rect 4869 144 4871 148
rect 4875 144 4877 148
rect 4881 144 4883 148
rect 4887 144 4889 148
rect 4893 144 4895 148
rect 4899 144 4901 148
rect 4905 144 4907 148
rect 4911 144 4913 148
rect 4917 144 4919 148
rect 4923 144 4925 148
rect 4929 144 4931 148
rect 4935 144 4937 148
rect 4941 144 4943 148
rect 4947 144 4949 148
rect 4953 144 4955 148
rect 4959 144 4961 148
rect 4965 144 4967 148
rect 4971 144 4973 148
rect 4977 144 4979 148
rect 4983 144 4985 148
rect 4989 144 4991 148
rect 4995 144 4998 148
rect 2 143 4998 144
<< nsubstratendiff >>
rect 4642 184 4680 187
rect 4642 180 4643 184
rect 4647 181 4675 184
rect 4647 180 4648 181
rect 4642 176 4648 180
rect 4674 180 4675 181
rect 4679 180 4680 184
rect 4642 172 4643 176
rect 4647 172 4648 176
rect 4642 168 4648 172
rect 4642 164 4643 168
rect 4647 164 4648 168
rect 4674 176 4680 180
rect 4674 172 4675 176
rect 4679 172 4680 176
rect 4674 168 4680 172
rect 4642 161 4648 164
rect 4674 164 4675 168
rect 4679 164 4680 168
rect 4674 161 4680 164
rect 4642 160 4680 161
rect 4642 156 4643 160
rect 4647 156 4655 160
rect 4659 156 4663 160
rect 4667 156 4675 160
rect 4679 156 4680 160
rect 4642 155 4680 156
rect 4698 184 4736 187
rect 4698 180 4699 184
rect 4703 181 4731 184
rect 4703 180 4704 181
rect 4698 176 4704 180
rect 4730 180 4731 181
rect 4735 180 4736 184
rect 4698 172 4699 176
rect 4703 172 4704 176
rect 4698 168 4704 172
rect 4698 164 4699 168
rect 4703 164 4704 168
rect 4730 176 4736 180
rect 4730 172 4731 176
rect 4735 172 4736 176
rect 4730 168 4736 172
rect 4698 161 4704 164
rect 4730 164 4731 168
rect 4735 164 4736 168
rect 4730 161 4736 164
rect 4698 160 4736 161
rect 4698 156 4699 160
rect 4703 156 4711 160
rect 4715 156 4719 160
rect 4723 156 4731 160
rect 4735 156 4736 160
rect 4698 155 4736 156
<< psubstratepcontact >>
rect 365 504 369 508
rect 365 498 369 502
rect 365 492 369 496
rect 365 486 369 490
rect 365 480 369 484
rect 365 474 369 478
rect 365 468 369 472
rect 365 462 369 466
rect 365 456 369 460
rect 365 450 369 454
rect 365 444 369 448
rect 365 438 369 442
rect 365 432 369 436
rect 365 426 369 430
rect 365 420 369 424
rect 365 414 369 418
rect 365 408 369 412
rect 365 402 369 406
rect 365 396 369 400
rect 365 390 369 394
rect 365 384 369 388
rect 365 378 369 382
rect 365 372 369 376
rect 365 366 369 370
rect 365 360 369 364
rect 365 354 369 358
rect 365 348 369 352
rect 365 342 369 346
rect 365 336 369 340
rect 365 330 369 334
rect 365 324 369 328
rect 365 318 369 322
rect 365 312 369 316
rect 365 306 369 310
rect 365 300 369 304
rect 365 294 369 298
rect 365 288 369 292
rect 365 282 369 286
rect 365 276 369 280
rect 365 270 369 274
rect 365 264 369 268
rect 365 258 369 262
rect 365 252 369 256
rect 365 246 369 250
rect 365 240 369 244
rect 365 234 369 238
rect 365 228 369 232
rect 365 222 369 226
rect 365 216 369 220
rect 365 210 369 214
rect 365 204 369 208
rect 365 198 369 202
rect 365 192 369 196
rect 365 186 369 190
rect 365 180 369 184
rect 365 174 369 178
rect 365 168 369 172
rect 365 162 369 166
rect 365 156 369 160
rect 365 150 369 154
rect 839 504 843 508
rect 839 498 843 502
rect 839 492 843 496
rect 839 486 843 490
rect 839 480 843 484
rect 839 474 843 478
rect 839 468 843 472
rect 839 462 843 466
rect 839 456 843 460
rect 839 450 843 454
rect 839 444 843 448
rect 839 438 843 442
rect 839 432 843 436
rect 839 426 843 430
rect 839 420 843 424
rect 839 414 843 418
rect 839 408 843 412
rect 839 402 843 406
rect 839 396 843 400
rect 839 390 843 394
rect 839 384 843 388
rect 839 378 843 382
rect 839 372 843 376
rect 839 366 843 370
rect 839 360 843 364
rect 839 354 843 358
rect 839 348 843 352
rect 839 342 843 346
rect 839 336 843 340
rect 839 330 843 334
rect 839 324 843 328
rect 839 318 843 322
rect 839 312 843 316
rect 839 306 843 310
rect 839 300 843 304
rect 839 294 843 298
rect 839 288 843 292
rect 839 282 843 286
rect 839 276 843 280
rect 839 270 843 274
rect 839 264 843 268
rect 839 258 843 262
rect 839 252 843 256
rect 839 246 843 250
rect 839 240 843 244
rect 839 234 843 238
rect 839 228 843 232
rect 839 222 843 226
rect 839 216 843 220
rect 839 210 843 214
rect 839 204 843 208
rect 839 198 843 202
rect 839 192 843 196
rect 839 186 843 190
rect 839 180 843 184
rect 839 174 843 178
rect 839 168 843 172
rect 839 162 843 166
rect 839 156 843 160
rect 839 150 843 154
rect 1313 504 1317 508
rect 1313 498 1317 502
rect 1313 492 1317 496
rect 1313 486 1317 490
rect 1313 480 1317 484
rect 1313 474 1317 478
rect 1313 468 1317 472
rect 1313 462 1317 466
rect 1313 456 1317 460
rect 1313 450 1317 454
rect 1313 444 1317 448
rect 1313 438 1317 442
rect 1313 432 1317 436
rect 1313 426 1317 430
rect 1313 420 1317 424
rect 1313 414 1317 418
rect 1313 408 1317 412
rect 1313 402 1317 406
rect 1313 396 1317 400
rect 1313 390 1317 394
rect 1313 384 1317 388
rect 1313 378 1317 382
rect 1313 372 1317 376
rect 1313 366 1317 370
rect 1313 360 1317 364
rect 1313 354 1317 358
rect 1313 348 1317 352
rect 1313 342 1317 346
rect 1313 336 1317 340
rect 1313 330 1317 334
rect 1313 324 1317 328
rect 1313 318 1317 322
rect 1313 312 1317 316
rect 1313 306 1317 310
rect 1313 300 1317 304
rect 1313 294 1317 298
rect 1313 288 1317 292
rect 1313 282 1317 286
rect 1313 276 1317 280
rect 1313 270 1317 274
rect 1313 264 1317 268
rect 1313 258 1317 262
rect 1313 252 1317 256
rect 1313 246 1317 250
rect 1313 240 1317 244
rect 1313 234 1317 238
rect 1313 228 1317 232
rect 1313 222 1317 226
rect 1313 216 1317 220
rect 1313 210 1317 214
rect 1313 204 1317 208
rect 1313 198 1317 202
rect 1313 192 1317 196
rect 1313 186 1317 190
rect 1313 180 1317 184
rect 1313 174 1317 178
rect 1313 168 1317 172
rect 1313 162 1317 166
rect 1313 156 1317 160
rect 1313 150 1317 154
rect 1787 504 1791 508
rect 1787 498 1791 502
rect 1787 492 1791 496
rect 1787 486 1791 490
rect 1787 480 1791 484
rect 1787 474 1791 478
rect 1787 468 1791 472
rect 1787 462 1791 466
rect 1787 456 1791 460
rect 1787 450 1791 454
rect 1787 444 1791 448
rect 1787 438 1791 442
rect 1787 432 1791 436
rect 1787 426 1791 430
rect 1787 420 1791 424
rect 1787 414 1791 418
rect 1787 408 1791 412
rect 1787 402 1791 406
rect 1787 396 1791 400
rect 1787 390 1791 394
rect 1787 384 1791 388
rect 1787 378 1791 382
rect 1787 372 1791 376
rect 1787 366 1791 370
rect 1787 360 1791 364
rect 1787 354 1791 358
rect 1787 348 1791 352
rect 1787 342 1791 346
rect 1787 336 1791 340
rect 1787 330 1791 334
rect 1787 324 1791 328
rect 1787 318 1791 322
rect 1787 312 1791 316
rect 1787 306 1791 310
rect 1787 300 1791 304
rect 1787 294 1791 298
rect 1787 288 1791 292
rect 1787 282 1791 286
rect 1787 276 1791 280
rect 1787 270 1791 274
rect 1787 264 1791 268
rect 1787 258 1791 262
rect 1787 252 1791 256
rect 1787 246 1791 250
rect 1787 240 1791 244
rect 1787 234 1791 238
rect 1787 228 1791 232
rect 1787 222 1791 226
rect 1787 216 1791 220
rect 1787 210 1791 214
rect 1787 204 1791 208
rect 1787 198 1791 202
rect 1787 192 1791 196
rect 1787 186 1791 190
rect 1787 180 1791 184
rect 1787 174 1791 178
rect 1787 168 1791 172
rect 1787 162 1791 166
rect 1787 156 1791 160
rect 1787 150 1791 154
rect 2261 504 2265 508
rect 2261 498 2265 502
rect 2261 492 2265 496
rect 2261 486 2265 490
rect 2261 480 2265 484
rect 2261 474 2265 478
rect 2261 468 2265 472
rect 2261 462 2265 466
rect 2261 456 2265 460
rect 2261 450 2265 454
rect 2261 444 2265 448
rect 2261 438 2265 442
rect 2261 432 2265 436
rect 2261 426 2265 430
rect 2261 420 2265 424
rect 2261 414 2265 418
rect 2261 408 2265 412
rect 2261 402 2265 406
rect 2261 396 2265 400
rect 2261 390 2265 394
rect 2261 384 2265 388
rect 2261 378 2265 382
rect 2261 372 2265 376
rect 2261 366 2265 370
rect 2261 360 2265 364
rect 2261 354 2265 358
rect 2261 348 2265 352
rect 2261 342 2265 346
rect 2261 336 2265 340
rect 2261 330 2265 334
rect 2261 324 2265 328
rect 2261 318 2265 322
rect 2261 312 2265 316
rect 2261 306 2265 310
rect 2261 300 2265 304
rect 2261 294 2265 298
rect 2261 288 2265 292
rect 2261 282 2265 286
rect 2261 276 2265 280
rect 2261 270 2265 274
rect 2261 264 2265 268
rect 2261 258 2265 262
rect 2261 252 2265 256
rect 2261 246 2265 250
rect 2261 240 2265 244
rect 2261 234 2265 238
rect 2261 228 2265 232
rect 2261 222 2265 226
rect 2261 216 2265 220
rect 2261 210 2265 214
rect 2261 204 2265 208
rect 2261 198 2265 202
rect 2261 192 2265 196
rect 2261 186 2265 190
rect 2261 180 2265 184
rect 2261 174 2265 178
rect 2261 168 2265 172
rect 2261 162 2265 166
rect 2261 156 2265 160
rect 2261 150 2265 154
rect 2735 504 2739 508
rect 2735 498 2739 502
rect 2735 492 2739 496
rect 2735 486 2739 490
rect 2735 480 2739 484
rect 2735 474 2739 478
rect 2735 468 2739 472
rect 2735 462 2739 466
rect 2735 456 2739 460
rect 2735 450 2739 454
rect 2735 444 2739 448
rect 2735 438 2739 442
rect 2735 432 2739 436
rect 2735 426 2739 430
rect 2735 420 2739 424
rect 2735 414 2739 418
rect 2735 408 2739 412
rect 2735 402 2739 406
rect 2735 396 2739 400
rect 2735 390 2739 394
rect 2735 384 2739 388
rect 2735 378 2739 382
rect 2735 372 2739 376
rect 2735 366 2739 370
rect 2735 360 2739 364
rect 2735 354 2739 358
rect 2735 348 2739 352
rect 2735 342 2739 346
rect 2735 336 2739 340
rect 2735 330 2739 334
rect 2735 324 2739 328
rect 2735 318 2739 322
rect 2735 312 2739 316
rect 2735 306 2739 310
rect 2735 300 2739 304
rect 2735 294 2739 298
rect 2735 288 2739 292
rect 2735 282 2739 286
rect 2735 276 2739 280
rect 2735 270 2739 274
rect 2735 264 2739 268
rect 2735 258 2739 262
rect 2735 252 2739 256
rect 2735 246 2739 250
rect 2735 240 2739 244
rect 2735 234 2739 238
rect 2735 228 2739 232
rect 2735 222 2739 226
rect 2735 216 2739 220
rect 2735 210 2739 214
rect 2735 204 2739 208
rect 2735 198 2739 202
rect 2735 192 2739 196
rect 2735 186 2739 190
rect 2735 180 2739 184
rect 2735 174 2739 178
rect 2735 168 2739 172
rect 2735 162 2739 166
rect 2735 156 2739 160
rect 2735 150 2739 154
rect 3209 504 3213 508
rect 3209 498 3213 502
rect 3209 492 3213 496
rect 3209 486 3213 490
rect 3209 480 3213 484
rect 3209 474 3213 478
rect 3209 468 3213 472
rect 3209 462 3213 466
rect 3209 456 3213 460
rect 3209 450 3213 454
rect 3209 444 3213 448
rect 3209 438 3213 442
rect 3209 432 3213 436
rect 3209 426 3213 430
rect 3209 420 3213 424
rect 3209 414 3213 418
rect 3209 408 3213 412
rect 3209 402 3213 406
rect 3209 396 3213 400
rect 3209 390 3213 394
rect 3209 384 3213 388
rect 3209 378 3213 382
rect 3209 372 3213 376
rect 3209 366 3213 370
rect 3209 360 3213 364
rect 3209 354 3213 358
rect 3209 348 3213 352
rect 3209 342 3213 346
rect 3209 336 3213 340
rect 3209 330 3213 334
rect 3209 324 3213 328
rect 3209 318 3213 322
rect 3209 312 3213 316
rect 3209 306 3213 310
rect 3209 300 3213 304
rect 3209 294 3213 298
rect 3209 288 3213 292
rect 3209 282 3213 286
rect 3209 276 3213 280
rect 3209 270 3213 274
rect 3209 264 3213 268
rect 3209 258 3213 262
rect 3209 252 3213 256
rect 3209 246 3213 250
rect 3209 240 3213 244
rect 3209 234 3213 238
rect 3209 228 3213 232
rect 3209 222 3213 226
rect 3209 216 3213 220
rect 3209 210 3213 214
rect 3209 204 3213 208
rect 3209 198 3213 202
rect 3209 192 3213 196
rect 3209 186 3213 190
rect 3209 180 3213 184
rect 3209 174 3213 178
rect 3209 168 3213 172
rect 3209 162 3213 166
rect 3209 156 3213 160
rect 3209 150 3213 154
rect 3683 504 3687 508
rect 3683 498 3687 502
rect 3683 492 3687 496
rect 3683 486 3687 490
rect 3683 480 3687 484
rect 3683 474 3687 478
rect 3683 468 3687 472
rect 3683 462 3687 466
rect 3683 456 3687 460
rect 3683 450 3687 454
rect 3683 444 3687 448
rect 3683 438 3687 442
rect 3683 432 3687 436
rect 3683 426 3687 430
rect 3683 420 3687 424
rect 3683 414 3687 418
rect 3683 408 3687 412
rect 3683 402 3687 406
rect 3683 396 3687 400
rect 3683 390 3687 394
rect 3683 384 3687 388
rect 3683 378 3687 382
rect 3683 372 3687 376
rect 3683 366 3687 370
rect 3683 360 3687 364
rect 3683 354 3687 358
rect 3683 348 3687 352
rect 3683 342 3687 346
rect 3683 336 3687 340
rect 3683 330 3687 334
rect 3683 324 3687 328
rect 3683 318 3687 322
rect 3683 312 3687 316
rect 3683 306 3687 310
rect 3683 300 3687 304
rect 3683 294 3687 298
rect 3683 288 3687 292
rect 3683 282 3687 286
rect 3683 276 3687 280
rect 3683 270 3687 274
rect 3683 264 3687 268
rect 3683 258 3687 262
rect 3683 252 3687 256
rect 3683 246 3687 250
rect 3683 240 3687 244
rect 3683 234 3687 238
rect 3683 228 3687 232
rect 3683 222 3687 226
rect 3683 216 3687 220
rect 3683 210 3687 214
rect 3683 204 3687 208
rect 3683 198 3687 202
rect 3683 192 3687 196
rect 3683 186 3687 190
rect 3683 180 3687 184
rect 3683 174 3687 178
rect 3683 168 3687 172
rect 3683 162 3687 166
rect 3683 156 3687 160
rect 3683 150 3687 154
rect 4157 504 4161 508
rect 4157 498 4161 502
rect 4157 492 4161 496
rect 4157 486 4161 490
rect 4157 480 4161 484
rect 4157 474 4161 478
rect 4157 468 4161 472
rect 4157 462 4161 466
rect 4157 456 4161 460
rect 4157 450 4161 454
rect 4157 444 4161 448
rect 4157 438 4161 442
rect 4157 432 4161 436
rect 4157 426 4161 430
rect 4157 420 4161 424
rect 4157 414 4161 418
rect 4157 408 4161 412
rect 4157 402 4161 406
rect 4157 396 4161 400
rect 4157 390 4161 394
rect 4157 384 4161 388
rect 4157 378 4161 382
rect 4157 372 4161 376
rect 4157 366 4161 370
rect 4157 360 4161 364
rect 4157 354 4161 358
rect 4157 348 4161 352
rect 4157 342 4161 346
rect 4157 336 4161 340
rect 4157 330 4161 334
rect 4157 324 4161 328
rect 4157 318 4161 322
rect 4157 312 4161 316
rect 4157 306 4161 310
rect 4157 300 4161 304
rect 4157 294 4161 298
rect 4157 288 4161 292
rect 4157 282 4161 286
rect 4157 276 4161 280
rect 4157 270 4161 274
rect 4157 264 4161 268
rect 4157 258 4161 262
rect 4157 252 4161 256
rect 4157 246 4161 250
rect 4157 240 4161 244
rect 4157 234 4161 238
rect 4157 228 4161 232
rect 4157 222 4161 226
rect 4157 216 4161 220
rect 4157 210 4161 214
rect 4157 204 4161 208
rect 4157 198 4161 202
rect 4157 192 4161 196
rect 4157 186 4161 190
rect 4157 180 4161 184
rect 4157 174 4161 178
rect 4157 168 4161 172
rect 4157 162 4161 166
rect 4157 156 4161 160
rect 4157 150 4161 154
rect 4631 504 4635 508
rect 4631 498 4635 502
rect 4631 492 4635 496
rect 4631 486 4635 490
rect 4631 480 4635 484
rect 4631 474 4635 478
rect 4631 468 4635 472
rect 4631 462 4635 466
rect 4631 456 4635 460
rect 4631 450 4635 454
rect 4631 444 4635 448
rect 4631 438 4635 442
rect 4631 432 4635 436
rect 4631 426 4635 430
rect 4631 420 4635 424
rect 4631 414 4635 418
rect 4631 408 4635 412
rect 4631 402 4635 406
rect 4631 396 4635 400
rect 4631 390 4635 394
rect 4631 384 4635 388
rect 4631 378 4635 382
rect 4631 372 4635 376
rect 4631 366 4635 370
rect 4631 360 4635 364
rect 4631 354 4635 358
rect 4631 348 4635 352
rect 4631 342 4635 346
rect 4631 336 4635 340
rect 4631 330 4635 334
rect 4631 324 4635 328
rect 4631 318 4635 322
rect 4631 312 4635 316
rect 4631 306 4635 310
rect 4631 300 4635 304
rect 4631 294 4635 298
rect 4631 288 4635 292
rect 4631 282 4635 286
rect 4631 276 4635 280
rect 4631 270 4635 274
rect 4631 264 4635 268
rect 4631 258 4635 262
rect 4631 252 4635 256
rect 4631 246 4635 250
rect 4631 240 4635 244
rect 4631 234 4635 238
rect 4631 228 4635 232
rect 4631 222 4635 226
rect 4631 216 4635 220
rect 4631 210 4635 214
rect 4631 204 4635 208
rect 4631 198 4635 202
rect 4631 192 4635 196
rect 4631 186 4635 190
rect 4631 180 4635 184
rect 4631 174 4635 178
rect 4631 168 4635 172
rect 4631 162 4635 166
rect 4631 156 4635 160
rect 4687 182 4691 186
rect 4687 176 4691 180
rect 4687 170 4691 174
rect 4687 164 4691 168
rect 4687 158 4691 162
rect 4631 150 4635 154
rect 4687 152 4691 156
rect 4743 182 4747 186
rect 4743 176 4747 180
rect 4743 170 4747 174
rect 4743 164 4747 168
rect 4743 158 4747 162
rect 4743 152 4747 156
rect 4769 182 4773 186
rect 4769 176 4773 180
rect 4769 170 4773 174
rect 4769 164 4773 168
rect 4769 158 4773 162
rect 4769 152 4773 156
rect 4795 182 4799 186
rect 4795 176 4799 180
rect 4795 170 4799 174
rect 4795 164 4799 168
rect 4795 158 4799 162
rect 4795 152 4799 156
rect 5 144 9 148
rect 11 144 15 148
rect 17 144 21 148
rect 23 144 27 148
rect 29 144 33 148
rect 35 144 39 148
rect 41 144 45 148
rect 47 144 51 148
rect 53 144 57 148
rect 59 144 63 148
rect 65 144 69 148
rect 71 144 75 148
rect 77 144 81 148
rect 83 144 87 148
rect 89 144 93 148
rect 95 144 99 148
rect 101 144 105 148
rect 107 144 111 148
rect 113 144 117 148
rect 119 144 123 148
rect 125 144 129 148
rect 131 144 135 148
rect 137 144 141 148
rect 143 144 147 148
rect 149 144 153 148
rect 155 144 159 148
rect 161 144 165 148
rect 167 144 171 148
rect 173 144 177 148
rect 179 144 183 148
rect 185 144 189 148
rect 191 144 195 148
rect 197 144 201 148
rect 203 144 207 148
rect 209 144 213 148
rect 215 144 219 148
rect 221 144 225 148
rect 227 144 231 148
rect 233 144 237 148
rect 239 144 243 148
rect 245 144 249 148
rect 251 144 255 148
rect 257 144 261 148
rect 263 144 267 148
rect 269 144 273 148
rect 275 144 279 148
rect 281 144 285 148
rect 287 144 291 148
rect 293 144 297 148
rect 299 144 303 148
rect 305 144 309 148
rect 311 144 315 148
rect 317 144 321 148
rect 323 144 327 148
rect 329 144 333 148
rect 335 144 339 148
rect 341 144 345 148
rect 347 144 351 148
rect 353 144 357 148
rect 359 144 363 148
rect 365 144 369 148
rect 371 144 375 148
rect 377 144 381 148
rect 383 144 387 148
rect 389 144 393 148
rect 395 144 399 148
rect 401 144 405 148
rect 407 144 411 148
rect 413 144 417 148
rect 419 144 423 148
rect 425 144 429 148
rect 431 144 435 148
rect 437 144 441 148
rect 443 144 447 148
rect 449 144 453 148
rect 455 144 459 148
rect 461 144 465 148
rect 467 144 471 148
rect 473 144 477 148
rect 479 144 483 148
rect 485 144 489 148
rect 491 144 495 148
rect 497 144 501 148
rect 503 144 507 148
rect 509 144 513 148
rect 515 144 519 148
rect 521 144 525 148
rect 527 144 531 148
rect 533 144 537 148
rect 539 144 543 148
rect 545 144 549 148
rect 551 144 555 148
rect 557 144 561 148
rect 563 144 567 148
rect 569 144 573 148
rect 575 144 579 148
rect 581 144 585 148
rect 587 144 591 148
rect 617 144 621 148
rect 623 144 627 148
rect 629 144 633 148
rect 635 144 639 148
rect 641 144 645 148
rect 647 144 651 148
rect 653 144 657 148
rect 659 144 663 148
rect 665 144 669 148
rect 671 144 675 148
rect 677 144 681 148
rect 683 144 687 148
rect 689 144 693 148
rect 695 144 699 148
rect 701 144 705 148
rect 707 144 711 148
rect 713 144 717 148
rect 719 144 723 148
rect 725 144 729 148
rect 731 144 735 148
rect 737 144 741 148
rect 743 144 747 148
rect 749 144 753 148
rect 755 144 759 148
rect 761 144 765 148
rect 767 144 771 148
rect 773 144 777 148
rect 779 144 783 148
rect 785 144 789 148
rect 791 144 795 148
rect 797 144 801 148
rect 803 144 807 148
rect 809 144 813 148
rect 815 144 819 148
rect 821 144 825 148
rect 827 144 831 148
rect 833 144 837 148
rect 839 144 843 148
rect 845 144 849 148
rect 851 144 855 148
rect 857 144 861 148
rect 863 144 867 148
rect 869 144 873 148
rect 875 144 879 148
rect 881 144 885 148
rect 887 144 891 148
rect 893 144 897 148
rect 899 144 903 148
rect 905 144 909 148
rect 911 144 915 148
rect 917 144 921 148
rect 923 144 927 148
rect 929 144 933 148
rect 935 144 939 148
rect 941 144 945 148
rect 947 144 951 148
rect 953 144 957 148
rect 959 144 963 148
rect 965 144 969 148
rect 971 144 975 148
rect 977 144 981 148
rect 983 144 987 148
rect 989 144 993 148
rect 995 144 999 148
rect 1001 144 1005 148
rect 1007 144 1011 148
rect 1013 144 1017 148
rect 1019 144 1023 148
rect 1025 144 1029 148
rect 1031 144 1035 148
rect 1037 144 1041 148
rect 1043 144 1047 148
rect 1049 144 1053 148
rect 1055 144 1059 148
rect 1061 144 1065 148
rect 1091 144 1095 148
rect 1097 144 1101 148
rect 1103 144 1107 148
rect 1109 144 1113 148
rect 1115 144 1119 148
rect 1121 144 1125 148
rect 1127 144 1131 148
rect 1133 144 1137 148
rect 1139 144 1143 148
rect 1145 144 1149 148
rect 1151 144 1155 148
rect 1157 144 1161 148
rect 1163 144 1167 148
rect 1169 144 1173 148
rect 1175 144 1179 148
rect 1181 144 1185 148
rect 1187 144 1191 148
rect 1193 144 1197 148
rect 1199 144 1203 148
rect 1205 144 1209 148
rect 1211 144 1215 148
rect 1217 144 1221 148
rect 1223 144 1227 148
rect 1229 144 1233 148
rect 1235 144 1239 148
rect 1241 144 1245 148
rect 1247 144 1251 148
rect 1253 144 1257 148
rect 1259 144 1263 148
rect 1265 144 1269 148
rect 1271 144 1275 148
rect 1277 144 1281 148
rect 1283 144 1287 148
rect 1289 144 1293 148
rect 1295 144 1299 148
rect 1301 144 1305 148
rect 1307 144 1311 148
rect 1313 144 1317 148
rect 1319 144 1323 148
rect 1325 144 1329 148
rect 1331 144 1335 148
rect 1337 144 1341 148
rect 1343 144 1347 148
rect 1349 144 1353 148
rect 1355 144 1359 148
rect 1361 144 1365 148
rect 1367 144 1371 148
rect 1373 144 1377 148
rect 1379 144 1383 148
rect 1385 144 1389 148
rect 1391 144 1395 148
rect 1397 144 1401 148
rect 1403 144 1407 148
rect 1409 144 1413 148
rect 1415 144 1419 148
rect 1421 144 1425 148
rect 1427 144 1431 148
rect 1433 144 1437 148
rect 1439 144 1443 148
rect 1445 144 1449 148
rect 1451 144 1455 148
rect 1457 144 1461 148
rect 1463 144 1467 148
rect 1469 144 1473 148
rect 1475 144 1479 148
rect 1481 144 1485 148
rect 1487 144 1491 148
rect 1493 144 1497 148
rect 1499 144 1503 148
rect 1505 144 1509 148
rect 1511 144 1515 148
rect 1517 144 1521 148
rect 1523 144 1527 148
rect 1529 144 1533 148
rect 1535 144 1539 148
rect 1565 144 1569 148
rect 1571 144 1575 148
rect 1577 144 1581 148
rect 1583 144 1587 148
rect 1589 144 1593 148
rect 1595 144 1599 148
rect 1601 144 1605 148
rect 1607 144 1611 148
rect 1613 144 1617 148
rect 1619 144 1623 148
rect 1625 144 1629 148
rect 1631 144 1635 148
rect 1637 144 1641 148
rect 1643 144 1647 148
rect 1649 144 1653 148
rect 1655 144 1659 148
rect 1661 144 1665 148
rect 1667 144 1671 148
rect 1673 144 1677 148
rect 1679 144 1683 148
rect 1685 144 1689 148
rect 1691 144 1695 148
rect 1697 144 1701 148
rect 1703 144 1707 148
rect 1709 144 1713 148
rect 1715 144 1719 148
rect 1721 144 1725 148
rect 1727 144 1731 148
rect 1733 144 1737 148
rect 1739 144 1743 148
rect 1745 144 1749 148
rect 1751 144 1755 148
rect 1757 144 1761 148
rect 1763 144 1767 148
rect 1769 144 1773 148
rect 1775 144 1779 148
rect 1781 144 1785 148
rect 1787 144 1791 148
rect 1793 144 1797 148
rect 1799 144 1803 148
rect 1805 144 1809 148
rect 1811 144 1815 148
rect 1817 144 1821 148
rect 1823 144 1827 148
rect 1829 144 1833 148
rect 1835 144 1839 148
rect 1841 144 1845 148
rect 1847 144 1851 148
rect 1853 144 1857 148
rect 1859 144 1863 148
rect 1865 144 1869 148
rect 1871 144 1875 148
rect 1877 144 1881 148
rect 1883 144 1887 148
rect 1889 144 1893 148
rect 1895 144 1899 148
rect 1901 144 1905 148
rect 1907 144 1911 148
rect 1913 144 1917 148
rect 1919 144 1923 148
rect 1925 144 1929 148
rect 1931 144 1935 148
rect 1937 144 1941 148
rect 1943 144 1947 148
rect 1949 144 1953 148
rect 1955 144 1959 148
rect 1961 144 1965 148
rect 1967 144 1971 148
rect 1973 144 1977 148
rect 1979 144 1983 148
rect 1985 144 1989 148
rect 1991 144 1995 148
rect 1997 144 2001 148
rect 2003 144 2007 148
rect 2009 144 2013 148
rect 2039 144 2043 148
rect 2045 144 2049 148
rect 2051 144 2055 148
rect 2057 144 2061 148
rect 2063 144 2067 148
rect 2069 144 2073 148
rect 2075 144 2079 148
rect 2081 144 2085 148
rect 2087 144 2091 148
rect 2093 144 2097 148
rect 2099 144 2103 148
rect 2105 144 2109 148
rect 2111 144 2115 148
rect 2117 144 2121 148
rect 2123 144 2127 148
rect 2129 144 2133 148
rect 2135 144 2139 148
rect 2141 144 2145 148
rect 2147 144 2151 148
rect 2153 144 2157 148
rect 2159 144 2163 148
rect 2165 144 2169 148
rect 2171 144 2175 148
rect 2177 144 2181 148
rect 2183 144 2187 148
rect 2189 144 2193 148
rect 2195 144 2199 148
rect 2201 144 2205 148
rect 2207 144 2211 148
rect 2213 144 2217 148
rect 2219 144 2223 148
rect 2225 144 2229 148
rect 2231 144 2235 148
rect 2237 144 2241 148
rect 2243 144 2247 148
rect 2249 144 2253 148
rect 2255 144 2259 148
rect 2261 144 2265 148
rect 2267 144 2271 148
rect 2273 144 2277 148
rect 2279 144 2283 148
rect 2285 144 2289 148
rect 2291 144 2295 148
rect 2297 144 2301 148
rect 2303 144 2307 148
rect 2309 144 2313 148
rect 2315 144 2319 148
rect 2321 144 2325 148
rect 2327 144 2331 148
rect 2333 144 2337 148
rect 2339 144 2343 148
rect 2345 144 2349 148
rect 2351 144 2355 148
rect 2357 144 2361 148
rect 2363 144 2367 148
rect 2369 144 2373 148
rect 2375 144 2379 148
rect 2381 144 2385 148
rect 2387 144 2391 148
rect 2393 144 2397 148
rect 2399 144 2403 148
rect 2405 144 2409 148
rect 2411 144 2415 148
rect 2417 144 2421 148
rect 2423 144 2427 148
rect 2429 144 2433 148
rect 2435 144 2439 148
rect 2441 144 2445 148
rect 2447 144 2451 148
rect 2453 144 2457 148
rect 2459 144 2463 148
rect 2465 144 2469 148
rect 2471 144 2475 148
rect 2477 144 2481 148
rect 2483 144 2487 148
rect 2513 144 2517 148
rect 2519 144 2523 148
rect 2525 144 2529 148
rect 2531 144 2535 148
rect 2537 144 2541 148
rect 2543 144 2547 148
rect 2549 144 2553 148
rect 2555 144 2559 148
rect 2561 144 2565 148
rect 2567 144 2571 148
rect 2573 144 2577 148
rect 2579 144 2583 148
rect 2585 144 2589 148
rect 2591 144 2595 148
rect 2597 144 2601 148
rect 2603 144 2607 148
rect 2609 144 2613 148
rect 2615 144 2619 148
rect 2621 144 2625 148
rect 2627 144 2631 148
rect 2633 144 2637 148
rect 2639 144 2643 148
rect 2645 144 2649 148
rect 2651 144 2655 148
rect 2657 144 2661 148
rect 2663 144 2667 148
rect 2669 144 2673 148
rect 2675 144 2679 148
rect 2681 144 2685 148
rect 2687 144 2691 148
rect 2693 144 2697 148
rect 2699 144 2703 148
rect 2705 144 2709 148
rect 2711 144 2715 148
rect 2717 144 2721 148
rect 2723 144 2727 148
rect 2729 144 2733 148
rect 2735 144 2739 148
rect 2741 144 2745 148
rect 2747 144 2751 148
rect 2753 144 2757 148
rect 2759 144 2763 148
rect 2765 144 2769 148
rect 2771 144 2775 148
rect 2777 144 2781 148
rect 2783 144 2787 148
rect 2789 144 2793 148
rect 2795 144 2799 148
rect 2801 144 2805 148
rect 2807 144 2811 148
rect 2813 144 2817 148
rect 2819 144 2823 148
rect 2825 144 2829 148
rect 2831 144 2835 148
rect 2837 144 2841 148
rect 2843 144 2847 148
rect 2849 144 2853 148
rect 2855 144 2859 148
rect 2861 144 2865 148
rect 2867 144 2871 148
rect 2873 144 2877 148
rect 2879 144 2883 148
rect 2885 144 2889 148
rect 2891 144 2895 148
rect 2897 144 2901 148
rect 2903 144 2907 148
rect 2909 144 2913 148
rect 2915 144 2919 148
rect 2921 144 2925 148
rect 2927 144 2931 148
rect 2933 144 2937 148
rect 2939 144 2943 148
rect 2945 144 2949 148
rect 2951 144 2955 148
rect 2957 144 2961 148
rect 2987 144 2991 148
rect 2993 144 2997 148
rect 2999 144 3003 148
rect 3005 144 3009 148
rect 3011 144 3015 148
rect 3017 144 3021 148
rect 3023 144 3027 148
rect 3029 144 3033 148
rect 3035 144 3039 148
rect 3041 144 3045 148
rect 3047 144 3051 148
rect 3053 144 3057 148
rect 3059 144 3063 148
rect 3065 144 3069 148
rect 3071 144 3075 148
rect 3077 144 3081 148
rect 3083 144 3087 148
rect 3089 144 3093 148
rect 3095 144 3099 148
rect 3101 144 3105 148
rect 3107 144 3111 148
rect 3113 144 3117 148
rect 3119 144 3123 148
rect 3125 144 3129 148
rect 3131 144 3135 148
rect 3137 144 3141 148
rect 3143 144 3147 148
rect 3149 144 3153 148
rect 3155 144 3159 148
rect 3161 144 3165 148
rect 3167 144 3171 148
rect 3173 144 3177 148
rect 3179 144 3183 148
rect 3185 144 3189 148
rect 3191 144 3195 148
rect 3197 144 3201 148
rect 3203 144 3207 148
rect 3209 144 3213 148
rect 3215 144 3219 148
rect 3221 144 3225 148
rect 3227 144 3231 148
rect 3233 144 3237 148
rect 3239 144 3243 148
rect 3245 144 3249 148
rect 3251 144 3255 148
rect 3257 144 3261 148
rect 3263 144 3267 148
rect 3269 144 3273 148
rect 3275 144 3279 148
rect 3281 144 3285 148
rect 3287 144 3291 148
rect 3293 144 3297 148
rect 3299 144 3303 148
rect 3305 144 3309 148
rect 3311 144 3315 148
rect 3317 144 3321 148
rect 3323 144 3327 148
rect 3329 144 3333 148
rect 3335 144 3339 148
rect 3341 144 3345 148
rect 3347 144 3351 148
rect 3353 144 3357 148
rect 3359 144 3363 148
rect 3365 144 3369 148
rect 3371 144 3375 148
rect 3377 144 3381 148
rect 3383 144 3387 148
rect 3389 144 3393 148
rect 3395 144 3399 148
rect 3401 144 3405 148
rect 3407 144 3411 148
rect 3413 144 3417 148
rect 3419 144 3423 148
rect 3425 144 3429 148
rect 3431 144 3435 148
rect 3461 144 3465 148
rect 3467 144 3471 148
rect 3473 144 3477 148
rect 3479 144 3483 148
rect 3485 144 3489 148
rect 3491 144 3495 148
rect 3497 144 3501 148
rect 3503 144 3507 148
rect 3509 144 3513 148
rect 3515 144 3519 148
rect 3521 144 3525 148
rect 3527 144 3531 148
rect 3533 144 3537 148
rect 3539 144 3543 148
rect 3545 144 3549 148
rect 3551 144 3555 148
rect 3557 144 3561 148
rect 3563 144 3567 148
rect 3569 144 3573 148
rect 3575 144 3579 148
rect 3581 144 3585 148
rect 3587 144 3591 148
rect 3593 144 3597 148
rect 3599 144 3603 148
rect 3605 144 3609 148
rect 3611 144 3615 148
rect 3617 144 3621 148
rect 3623 144 3627 148
rect 3629 144 3633 148
rect 3635 144 3639 148
rect 3641 144 3645 148
rect 3647 144 3651 148
rect 3653 144 3657 148
rect 3659 144 3663 148
rect 3665 144 3669 148
rect 3671 144 3675 148
rect 3677 144 3681 148
rect 3683 144 3687 148
rect 3689 144 3693 148
rect 3695 144 3699 148
rect 3701 144 3705 148
rect 3707 144 3711 148
rect 3713 144 3717 148
rect 3719 144 3723 148
rect 3725 144 3729 148
rect 3731 144 3735 148
rect 3737 144 3741 148
rect 3743 144 3747 148
rect 3749 144 3753 148
rect 3755 144 3759 148
rect 3761 144 3765 148
rect 3767 144 3771 148
rect 3773 144 3777 148
rect 3779 144 3783 148
rect 3785 144 3789 148
rect 3791 144 3795 148
rect 3797 144 3801 148
rect 3803 144 3807 148
rect 3809 144 3813 148
rect 3815 144 3819 148
rect 3821 144 3825 148
rect 3827 144 3831 148
rect 3833 144 3837 148
rect 3839 144 3843 148
rect 3845 144 3849 148
rect 3851 144 3855 148
rect 3857 144 3861 148
rect 3863 144 3867 148
rect 3869 144 3873 148
rect 3875 144 3879 148
rect 3881 144 3885 148
rect 3887 144 3891 148
rect 3893 144 3897 148
rect 3899 144 3903 148
rect 3905 144 3909 148
rect 3935 144 3939 148
rect 3941 144 3945 148
rect 3947 144 3951 148
rect 3953 144 3957 148
rect 3959 144 3963 148
rect 3965 144 3969 148
rect 3971 144 3975 148
rect 3977 144 3981 148
rect 3983 144 3987 148
rect 3989 144 3993 148
rect 3995 144 3999 148
rect 4001 144 4005 148
rect 4007 144 4011 148
rect 4013 144 4017 148
rect 4019 144 4023 148
rect 4025 144 4029 148
rect 4031 144 4035 148
rect 4037 144 4041 148
rect 4043 144 4047 148
rect 4049 144 4053 148
rect 4055 144 4059 148
rect 4061 144 4065 148
rect 4067 144 4071 148
rect 4073 144 4077 148
rect 4079 144 4083 148
rect 4085 144 4089 148
rect 4091 144 4095 148
rect 4097 144 4101 148
rect 4103 144 4107 148
rect 4109 144 4113 148
rect 4115 144 4119 148
rect 4121 144 4125 148
rect 4127 144 4131 148
rect 4133 144 4137 148
rect 4139 144 4143 148
rect 4145 144 4149 148
rect 4151 144 4155 148
rect 4157 144 4161 148
rect 4163 144 4167 148
rect 4169 144 4173 148
rect 4175 144 4179 148
rect 4181 144 4185 148
rect 4187 144 4191 148
rect 4193 144 4197 148
rect 4199 144 4203 148
rect 4205 144 4209 148
rect 4211 144 4215 148
rect 4217 144 4221 148
rect 4223 144 4227 148
rect 4229 144 4233 148
rect 4235 144 4239 148
rect 4241 144 4245 148
rect 4247 144 4251 148
rect 4253 144 4257 148
rect 4259 144 4263 148
rect 4265 144 4269 148
rect 4271 144 4275 148
rect 4277 144 4281 148
rect 4283 144 4287 148
rect 4289 144 4293 148
rect 4295 144 4299 148
rect 4301 144 4305 148
rect 4307 144 4311 148
rect 4313 144 4317 148
rect 4319 144 4323 148
rect 4325 144 4329 148
rect 4331 144 4335 148
rect 4337 144 4341 148
rect 4343 144 4347 148
rect 4349 144 4353 148
rect 4355 144 4359 148
rect 4361 144 4365 148
rect 4367 144 4371 148
rect 4373 144 4377 148
rect 4379 144 4383 148
rect 4409 144 4413 148
rect 4415 144 4419 148
rect 4421 144 4425 148
rect 4427 144 4431 148
rect 4433 144 4437 148
rect 4439 144 4443 148
rect 4445 144 4449 148
rect 4451 144 4455 148
rect 4457 144 4461 148
rect 4463 144 4467 148
rect 4469 144 4473 148
rect 4475 144 4479 148
rect 4481 144 4485 148
rect 4487 144 4491 148
rect 4493 144 4497 148
rect 4499 144 4503 148
rect 4505 144 4509 148
rect 4511 144 4515 148
rect 4517 144 4521 148
rect 4523 144 4527 148
rect 4529 144 4533 148
rect 4535 144 4539 148
rect 4541 144 4545 148
rect 4547 144 4551 148
rect 4553 144 4557 148
rect 4559 144 4563 148
rect 4565 144 4569 148
rect 4571 144 4575 148
rect 4577 144 4581 148
rect 4583 144 4587 148
rect 4589 144 4593 148
rect 4595 144 4599 148
rect 4601 144 4605 148
rect 4607 144 4611 148
rect 4613 144 4617 148
rect 4619 144 4623 148
rect 4625 144 4629 148
rect 4631 144 4635 148
rect 4637 144 4641 148
rect 4643 144 4647 148
rect 4649 144 4653 148
rect 4655 144 4659 148
rect 4661 144 4665 148
rect 4667 144 4671 148
rect 4673 144 4677 148
rect 4679 144 4683 148
rect 4685 144 4689 148
rect 4691 144 4695 148
rect 4697 144 4701 148
rect 4703 144 4707 148
rect 4709 144 4713 148
rect 4715 144 4719 148
rect 4721 144 4725 148
rect 4727 144 4731 148
rect 4733 144 4737 148
rect 4739 144 4743 148
rect 4745 144 4749 148
rect 4751 144 4755 148
rect 4757 144 4761 148
rect 4763 144 4767 148
rect 4769 144 4773 148
rect 4775 144 4779 148
rect 4781 144 4785 148
rect 4787 144 4791 148
rect 4793 144 4797 148
rect 4799 144 4803 148
rect 4805 144 4809 148
rect 4811 144 4815 148
rect 4817 144 4821 148
rect 4823 144 4827 148
rect 4829 144 4833 148
rect 4835 144 4839 148
rect 4841 144 4845 148
rect 4847 144 4851 148
rect 4853 144 4857 148
rect 4859 144 4863 148
rect 4865 144 4869 148
rect 4871 144 4875 148
rect 4877 144 4881 148
rect 4883 144 4887 148
rect 4889 144 4893 148
rect 4895 144 4899 148
rect 4901 144 4905 148
rect 4907 144 4911 148
rect 4913 144 4917 148
rect 4919 144 4923 148
rect 4925 144 4929 148
rect 4931 144 4935 148
rect 4937 144 4941 148
rect 4943 144 4947 148
rect 4949 144 4953 148
rect 4955 144 4959 148
rect 4961 144 4965 148
rect 4967 144 4971 148
rect 4973 144 4977 148
rect 4979 144 4983 148
rect 4985 144 4989 148
rect 4991 144 4995 148
<< nsubstratencontact >>
rect 4643 180 4647 184
rect 4675 180 4679 184
rect 4643 172 4647 176
rect 4643 164 4647 168
rect 4675 172 4679 176
rect 4675 164 4679 168
rect 4643 156 4647 160
rect 4655 156 4659 160
rect 4663 156 4667 160
rect 4675 156 4679 160
rect 4699 180 4703 184
rect 4731 180 4735 184
rect 4699 172 4703 176
rect 4699 164 4703 168
rect 4731 172 4735 176
rect 4731 164 4735 168
rect 4699 156 4703 160
rect 4711 156 4715 160
rect 4719 156 4723 160
rect 4731 156 4735 160
<< polysilicon >>
rect 4642 499 4685 501
rect 4642 490 4669 499
rect 4683 490 4685 499
rect 4642 488 4685 490
rect 4642 222 4654 488
rect 4657 473 4684 485
rect 4657 222 4669 473
rect 4642 210 4669 222
rect 4672 228 4684 473
rect 4672 226 4685 228
rect 4672 212 4674 226
rect 4683 212 4685 226
rect 4672 210 4685 212
rect 4811 196 4824 198
rect 4970 197 4988 198
rect 4811 182 4813 196
rect 4822 182 4824 196
rect 4811 167 4824 182
rect 4827 196 4988 197
rect 4827 187 4972 196
rect 4986 187 4988 196
rect 4827 185 4988 187
rect 4827 182 4839 185
rect 4827 170 4988 182
rect 4976 167 4988 170
rect 4811 155 4988 167
rect 371 141 4629 142
rect 371 137 495 141
rect 499 137 501 141
rect 505 137 507 141
rect 511 137 513 141
rect 517 137 519 141
rect 523 137 525 141
rect 529 137 531 141
rect 535 137 673 141
rect 677 137 679 141
rect 683 137 685 141
rect 689 137 691 141
rect 695 137 697 141
rect 701 137 703 141
rect 707 137 709 141
rect 713 137 969 141
rect 973 137 975 141
rect 979 137 981 141
rect 985 137 987 141
rect 991 137 993 141
rect 997 137 999 141
rect 1003 137 1005 141
rect 1009 137 1147 141
rect 1151 137 1153 141
rect 1157 137 1159 141
rect 1163 137 1165 141
rect 1169 137 1171 141
rect 1175 137 1177 141
rect 1181 137 1183 141
rect 1187 137 1443 141
rect 1447 137 1449 141
rect 1453 137 1455 141
rect 1459 137 1461 141
rect 1465 137 1467 141
rect 1471 137 1473 141
rect 1477 137 1479 141
rect 1483 137 1621 141
rect 1625 137 1627 141
rect 1631 137 1633 141
rect 1637 137 1639 141
rect 1643 137 1645 141
rect 1649 137 1651 141
rect 1655 137 1657 141
rect 1661 137 1917 141
rect 1921 137 1923 141
rect 1927 137 1929 141
rect 1933 137 1935 141
rect 1939 137 1941 141
rect 1945 137 1947 141
rect 1951 137 1953 141
rect 1957 137 2095 141
rect 2099 137 2101 141
rect 2105 137 2107 141
rect 2111 137 2113 141
rect 2117 137 2119 141
rect 2123 137 2125 141
rect 2129 137 2131 141
rect 2135 137 2391 141
rect 2395 137 2397 141
rect 2401 137 2403 141
rect 2407 137 2409 141
rect 2413 137 2415 141
rect 2419 137 2421 141
rect 2425 137 2427 141
rect 2431 137 2569 141
rect 2573 137 2575 141
rect 2579 137 2581 141
rect 2585 137 2587 141
rect 2591 137 2593 141
rect 2597 137 2599 141
rect 2603 137 2605 141
rect 2609 137 2865 141
rect 2869 137 2871 141
rect 2875 137 2877 141
rect 2881 137 2883 141
rect 2887 137 2889 141
rect 2893 137 2895 141
rect 2899 137 2901 141
rect 2905 137 3043 141
rect 3047 137 3049 141
rect 3053 137 3055 141
rect 3059 137 3061 141
rect 3065 137 3067 141
rect 3071 137 3073 141
rect 3077 137 3079 141
rect 3083 137 3339 141
rect 3343 137 3345 141
rect 3349 137 3351 141
rect 3355 137 3357 141
rect 3361 137 3363 141
rect 3367 137 3369 141
rect 3373 137 3375 141
rect 3379 137 3517 141
rect 3521 137 3523 141
rect 3527 137 3529 141
rect 3533 137 3535 141
rect 3539 137 3541 141
rect 3545 137 3547 141
rect 3551 137 3553 141
rect 3557 137 3813 141
rect 3817 137 3819 141
rect 3823 137 3825 141
rect 3829 137 3831 141
rect 3835 137 3837 141
rect 3841 137 3843 141
rect 3847 137 3849 141
rect 3853 137 3991 141
rect 3995 137 3997 141
rect 4001 137 4003 141
rect 4007 137 4009 141
rect 4013 137 4015 141
rect 4019 137 4021 141
rect 4025 137 4027 141
rect 4031 137 4287 141
rect 4291 137 4293 141
rect 4297 137 4299 141
rect 4303 137 4305 141
rect 4309 137 4311 141
rect 4315 137 4317 141
rect 4321 137 4323 141
rect 4327 137 4465 141
rect 4469 137 4471 141
rect 4475 137 4477 141
rect 4481 137 4483 141
rect 4487 137 4489 141
rect 4493 137 4495 141
rect 4499 137 4501 141
rect 4505 137 4629 141
rect 371 12 4629 137
rect 371 8 673 12
rect 677 8 679 12
rect 683 8 685 12
rect 689 8 691 12
rect 695 8 697 12
rect 701 8 703 12
rect 707 8 709 12
rect 713 8 969 12
rect 973 8 975 12
rect 979 8 981 12
rect 985 8 987 12
rect 991 8 993 12
rect 997 8 999 12
rect 1003 8 1005 12
rect 1009 8 1147 12
rect 1151 8 1153 12
rect 1157 8 1159 12
rect 1163 8 1165 12
rect 1169 8 1171 12
rect 1175 8 1177 12
rect 1181 8 1183 12
rect 1187 8 1443 12
rect 1447 8 1449 12
rect 1453 8 1455 12
rect 1459 8 1461 12
rect 1465 8 1467 12
rect 1471 8 1473 12
rect 1477 8 1479 12
rect 1483 8 1621 12
rect 1625 8 1627 12
rect 1631 8 1633 12
rect 1637 8 1639 12
rect 1643 8 1645 12
rect 1649 8 1651 12
rect 1655 8 1657 12
rect 1661 8 1917 12
rect 1921 8 1923 12
rect 1927 8 1929 12
rect 1933 8 1935 12
rect 1939 8 1941 12
rect 1945 8 1947 12
rect 1951 8 1953 12
rect 1957 8 2095 12
rect 2099 8 2101 12
rect 2105 8 2107 12
rect 2111 8 2113 12
rect 2117 8 2119 12
rect 2123 8 2125 12
rect 2129 8 2131 12
rect 2135 8 2391 12
rect 2395 8 2397 12
rect 2401 8 2403 12
rect 2407 8 2409 12
rect 2413 8 2415 12
rect 2419 8 2421 12
rect 2425 8 2427 12
rect 2431 8 2569 12
rect 2573 8 2575 12
rect 2579 8 2581 12
rect 2585 8 2587 12
rect 2591 8 2593 12
rect 2597 8 2599 12
rect 2603 8 2605 12
rect 2609 8 2865 12
rect 2869 8 2871 12
rect 2875 8 2877 12
rect 2881 8 2883 12
rect 2887 8 2889 12
rect 2893 8 2895 12
rect 2899 8 2901 12
rect 2905 8 3043 12
rect 3047 8 3049 12
rect 3053 8 3055 12
rect 3059 8 3061 12
rect 3065 8 3067 12
rect 3071 8 3073 12
rect 3077 8 3079 12
rect 3083 8 3339 12
rect 3343 8 3345 12
rect 3349 8 3351 12
rect 3355 8 3357 12
rect 3361 8 3363 12
rect 3367 8 3369 12
rect 3373 8 3375 12
rect 3379 8 3517 12
rect 3521 8 3523 12
rect 3527 8 3529 12
rect 3533 8 3535 12
rect 3539 8 3541 12
rect 3545 8 3547 12
rect 3551 8 3553 12
rect 3557 8 3813 12
rect 3817 8 3819 12
rect 3823 8 3825 12
rect 3829 8 3831 12
rect 3835 8 3837 12
rect 3841 8 3843 12
rect 3847 8 3849 12
rect 3853 8 3991 12
rect 3995 8 3997 12
rect 4001 8 4003 12
rect 4007 8 4009 12
rect 4013 8 4015 12
rect 4019 8 4021 12
rect 4025 8 4027 12
rect 4031 8 4287 12
rect 4291 8 4293 12
rect 4297 8 4299 12
rect 4303 8 4305 12
rect 4309 8 4311 12
rect 4315 8 4317 12
rect 4321 8 4323 12
rect 4327 8 4629 12
rect 371 7 4629 8
<< polycontact >>
rect 4669 490 4683 499
rect 4674 212 4683 226
rect 4813 182 4822 196
rect 4972 187 4986 196
rect 495 137 499 141
rect 501 137 505 141
rect 507 137 511 141
rect 513 137 517 141
rect 519 137 523 141
rect 525 137 529 141
rect 531 137 535 141
rect 673 137 677 141
rect 679 137 683 141
rect 685 137 689 141
rect 691 137 695 141
rect 697 137 701 141
rect 703 137 707 141
rect 709 137 713 141
rect 969 137 973 141
rect 975 137 979 141
rect 981 137 985 141
rect 987 137 991 141
rect 993 137 997 141
rect 999 137 1003 141
rect 1005 137 1009 141
rect 1147 137 1151 141
rect 1153 137 1157 141
rect 1159 137 1163 141
rect 1165 137 1169 141
rect 1171 137 1175 141
rect 1177 137 1181 141
rect 1183 137 1187 141
rect 1443 137 1447 141
rect 1449 137 1453 141
rect 1455 137 1459 141
rect 1461 137 1465 141
rect 1467 137 1471 141
rect 1473 137 1477 141
rect 1479 137 1483 141
rect 1621 137 1625 141
rect 1627 137 1631 141
rect 1633 137 1637 141
rect 1639 137 1643 141
rect 1645 137 1649 141
rect 1651 137 1655 141
rect 1657 137 1661 141
rect 1917 137 1921 141
rect 1923 137 1927 141
rect 1929 137 1933 141
rect 1935 137 1939 141
rect 1941 137 1945 141
rect 1947 137 1951 141
rect 1953 137 1957 141
rect 2095 137 2099 141
rect 2101 137 2105 141
rect 2107 137 2111 141
rect 2113 137 2117 141
rect 2119 137 2123 141
rect 2125 137 2129 141
rect 2131 137 2135 141
rect 2391 137 2395 141
rect 2397 137 2401 141
rect 2403 137 2407 141
rect 2409 137 2413 141
rect 2415 137 2419 141
rect 2421 137 2425 141
rect 2427 137 2431 141
rect 2569 137 2573 141
rect 2575 137 2579 141
rect 2581 137 2585 141
rect 2587 137 2591 141
rect 2593 137 2597 141
rect 2599 137 2603 141
rect 2605 137 2609 141
rect 2865 137 2869 141
rect 2871 137 2875 141
rect 2877 137 2881 141
rect 2883 137 2887 141
rect 2889 137 2893 141
rect 2895 137 2899 141
rect 2901 137 2905 141
rect 3043 137 3047 141
rect 3049 137 3053 141
rect 3055 137 3059 141
rect 3061 137 3065 141
rect 3067 137 3071 141
rect 3073 137 3077 141
rect 3079 137 3083 141
rect 3339 137 3343 141
rect 3345 137 3349 141
rect 3351 137 3355 141
rect 3357 137 3361 141
rect 3363 137 3367 141
rect 3369 137 3373 141
rect 3375 137 3379 141
rect 3517 137 3521 141
rect 3523 137 3527 141
rect 3529 137 3533 141
rect 3535 137 3539 141
rect 3541 137 3545 141
rect 3547 137 3551 141
rect 3553 137 3557 141
rect 3813 137 3817 141
rect 3819 137 3823 141
rect 3825 137 3829 141
rect 3831 137 3835 141
rect 3837 137 3841 141
rect 3843 137 3847 141
rect 3849 137 3853 141
rect 3991 137 3995 141
rect 3997 137 4001 141
rect 4003 137 4007 141
rect 4009 137 4013 141
rect 4015 137 4019 141
rect 4021 137 4025 141
rect 4027 137 4031 141
rect 4287 137 4291 141
rect 4293 137 4297 141
rect 4299 137 4303 141
rect 4305 137 4309 141
rect 4311 137 4315 141
rect 4317 137 4321 141
rect 4323 137 4327 141
rect 4465 137 4469 141
rect 4471 137 4475 141
rect 4477 137 4481 141
rect 4483 137 4487 141
rect 4489 137 4493 141
rect 4495 137 4499 141
rect 4501 137 4505 141
rect 673 8 677 12
rect 679 8 683 12
rect 685 8 689 12
rect 691 8 695 12
rect 697 8 701 12
rect 703 8 707 12
rect 709 8 713 12
rect 969 8 973 12
rect 975 8 979 12
rect 981 8 985 12
rect 987 8 991 12
rect 993 8 997 12
rect 999 8 1003 12
rect 1005 8 1009 12
rect 1147 8 1151 12
rect 1153 8 1157 12
rect 1159 8 1163 12
rect 1165 8 1169 12
rect 1171 8 1175 12
rect 1177 8 1181 12
rect 1183 8 1187 12
rect 1443 8 1447 12
rect 1449 8 1453 12
rect 1455 8 1459 12
rect 1461 8 1465 12
rect 1467 8 1471 12
rect 1473 8 1477 12
rect 1479 8 1483 12
rect 1621 8 1625 12
rect 1627 8 1631 12
rect 1633 8 1637 12
rect 1639 8 1643 12
rect 1645 8 1649 12
rect 1651 8 1655 12
rect 1657 8 1661 12
rect 1917 8 1921 12
rect 1923 8 1927 12
rect 1929 8 1933 12
rect 1935 8 1939 12
rect 1941 8 1945 12
rect 1947 8 1951 12
rect 1953 8 1957 12
rect 2095 8 2099 12
rect 2101 8 2105 12
rect 2107 8 2111 12
rect 2113 8 2117 12
rect 2119 8 2123 12
rect 2125 8 2129 12
rect 2131 8 2135 12
rect 2391 8 2395 12
rect 2397 8 2401 12
rect 2403 8 2407 12
rect 2409 8 2413 12
rect 2415 8 2419 12
rect 2421 8 2425 12
rect 2427 8 2431 12
rect 2569 8 2573 12
rect 2575 8 2579 12
rect 2581 8 2585 12
rect 2587 8 2591 12
rect 2593 8 2597 12
rect 2599 8 2603 12
rect 2605 8 2609 12
rect 2865 8 2869 12
rect 2871 8 2875 12
rect 2877 8 2881 12
rect 2883 8 2887 12
rect 2889 8 2893 12
rect 2895 8 2899 12
rect 2901 8 2905 12
rect 3043 8 3047 12
rect 3049 8 3053 12
rect 3055 8 3059 12
rect 3061 8 3065 12
rect 3067 8 3071 12
rect 3073 8 3077 12
rect 3079 8 3083 12
rect 3339 8 3343 12
rect 3345 8 3349 12
rect 3351 8 3355 12
rect 3357 8 3361 12
rect 3363 8 3367 12
rect 3369 8 3373 12
rect 3375 8 3379 12
rect 3517 8 3521 12
rect 3523 8 3527 12
rect 3529 8 3533 12
rect 3535 8 3539 12
rect 3541 8 3545 12
rect 3547 8 3551 12
rect 3553 8 3557 12
rect 3813 8 3817 12
rect 3819 8 3823 12
rect 3825 8 3829 12
rect 3831 8 3835 12
rect 3837 8 3841 12
rect 3843 8 3847 12
rect 3849 8 3853 12
rect 3991 8 3995 12
rect 3997 8 4001 12
rect 4003 8 4007 12
rect 4009 8 4013 12
rect 4015 8 4019 12
rect 4021 8 4025 12
rect 4027 8 4031 12
rect 4287 8 4291 12
rect 4293 8 4297 12
rect 4299 8 4303 12
rect 4305 8 4309 12
rect 4311 8 4315 12
rect 4317 8 4321 12
rect 4323 8 4327 12
<< metal1 >>
rect 365 508 369 510
rect 365 502 369 504
rect 365 496 369 498
rect 365 490 369 492
rect 365 484 369 486
rect 365 478 369 480
rect 365 472 369 474
rect 365 466 369 468
rect 365 460 369 462
rect 365 454 369 456
rect 365 448 369 450
rect 365 442 369 444
rect 365 436 369 438
rect 365 430 369 432
rect 365 424 369 426
rect 365 418 369 420
rect 365 412 369 414
rect 365 406 369 408
rect 365 400 369 402
rect 365 394 369 396
rect 365 388 369 390
rect 365 382 369 384
rect 365 376 369 378
rect 365 370 369 372
rect 365 364 369 366
rect 365 358 369 360
rect 365 352 369 354
rect 365 346 369 348
rect 365 340 369 342
rect 365 334 369 336
rect 365 328 369 330
rect 365 322 369 324
rect 365 316 369 318
rect 365 310 369 312
rect 365 304 369 306
rect 365 298 369 300
rect 365 292 369 294
rect 365 286 369 288
rect 365 280 369 282
rect 365 274 369 276
rect 365 268 369 270
rect 365 262 369 264
rect 365 256 369 258
rect 365 250 369 252
rect 365 244 369 246
rect 365 238 369 240
rect 365 232 369 234
rect 365 226 369 228
rect 365 220 369 222
rect 365 214 369 216
rect 365 208 369 210
rect 365 202 369 204
rect 365 196 369 198
rect 365 190 369 192
rect 365 184 369 186
rect 365 178 369 180
rect 365 172 369 174
rect 365 166 369 168
rect 365 160 369 162
rect 365 154 369 156
rect 365 148 369 150
rect 839 508 843 510
rect 839 502 843 504
rect 839 496 843 498
rect 839 490 843 492
rect 839 484 843 486
rect 839 478 843 480
rect 839 472 843 474
rect 839 466 843 468
rect 839 460 843 462
rect 839 454 843 456
rect 839 448 843 450
rect 839 442 843 444
rect 839 436 843 438
rect 839 430 843 432
rect 839 424 843 426
rect 839 418 843 420
rect 839 412 843 414
rect 839 406 843 408
rect 839 400 843 402
rect 839 394 843 396
rect 839 388 843 390
rect 839 382 843 384
rect 839 376 843 378
rect 839 370 843 372
rect 839 364 843 366
rect 839 358 843 360
rect 839 352 843 354
rect 839 346 843 348
rect 839 340 843 342
rect 839 334 843 336
rect 839 328 843 330
rect 839 322 843 324
rect 839 316 843 318
rect 839 310 843 312
rect 839 304 843 306
rect 839 298 843 300
rect 839 292 843 294
rect 839 286 843 288
rect 839 280 843 282
rect 839 274 843 276
rect 839 268 843 270
rect 839 262 843 264
rect 839 256 843 258
rect 839 250 843 252
rect 839 244 843 246
rect 839 238 843 240
rect 839 232 843 234
rect 839 226 843 228
rect 839 220 843 222
rect 839 214 843 216
rect 839 208 843 210
rect 839 202 843 204
rect 839 196 843 198
rect 839 190 843 192
rect 839 184 843 186
rect 839 178 843 180
rect 839 172 843 174
rect 839 166 843 168
rect 839 160 843 162
rect 839 154 843 156
rect 839 148 843 150
rect 1313 508 1317 510
rect 1313 502 1317 504
rect 1313 496 1317 498
rect 1313 490 1317 492
rect 1313 484 1317 486
rect 1313 478 1317 480
rect 1313 472 1317 474
rect 1313 466 1317 468
rect 1313 460 1317 462
rect 1313 454 1317 456
rect 1313 448 1317 450
rect 1313 442 1317 444
rect 1313 436 1317 438
rect 1313 430 1317 432
rect 1313 424 1317 426
rect 1313 418 1317 420
rect 1313 412 1317 414
rect 1313 406 1317 408
rect 1313 400 1317 402
rect 1313 394 1317 396
rect 1313 388 1317 390
rect 1313 382 1317 384
rect 1313 376 1317 378
rect 1313 370 1317 372
rect 1313 364 1317 366
rect 1313 358 1317 360
rect 1313 352 1317 354
rect 1313 346 1317 348
rect 1313 340 1317 342
rect 1313 334 1317 336
rect 1313 328 1317 330
rect 1313 322 1317 324
rect 1313 316 1317 318
rect 1313 310 1317 312
rect 1313 304 1317 306
rect 1313 298 1317 300
rect 1313 292 1317 294
rect 1313 286 1317 288
rect 1313 280 1317 282
rect 1313 274 1317 276
rect 1313 268 1317 270
rect 1313 262 1317 264
rect 1313 256 1317 258
rect 1313 250 1317 252
rect 1313 244 1317 246
rect 1313 238 1317 240
rect 1313 232 1317 234
rect 1313 226 1317 228
rect 1313 220 1317 222
rect 1313 214 1317 216
rect 1313 208 1317 210
rect 1313 202 1317 204
rect 1313 196 1317 198
rect 1313 190 1317 192
rect 1313 184 1317 186
rect 1313 178 1317 180
rect 1313 172 1317 174
rect 1313 166 1317 168
rect 1313 160 1317 162
rect 1313 154 1317 156
rect 1313 148 1317 150
rect 1787 508 1791 510
rect 1787 502 1791 504
rect 1787 496 1791 498
rect 1787 490 1791 492
rect 1787 484 1791 486
rect 1787 478 1791 480
rect 1787 472 1791 474
rect 1787 466 1791 468
rect 1787 460 1791 462
rect 1787 454 1791 456
rect 1787 448 1791 450
rect 1787 442 1791 444
rect 1787 436 1791 438
rect 1787 430 1791 432
rect 1787 424 1791 426
rect 1787 418 1791 420
rect 1787 412 1791 414
rect 1787 406 1791 408
rect 1787 400 1791 402
rect 1787 394 1791 396
rect 1787 388 1791 390
rect 1787 382 1791 384
rect 1787 376 1791 378
rect 1787 370 1791 372
rect 1787 364 1791 366
rect 1787 358 1791 360
rect 1787 352 1791 354
rect 1787 346 1791 348
rect 1787 340 1791 342
rect 1787 334 1791 336
rect 1787 328 1791 330
rect 1787 322 1791 324
rect 1787 316 1791 318
rect 1787 310 1791 312
rect 1787 304 1791 306
rect 1787 298 1791 300
rect 1787 292 1791 294
rect 1787 286 1791 288
rect 1787 280 1791 282
rect 1787 274 1791 276
rect 1787 268 1791 270
rect 1787 262 1791 264
rect 1787 256 1791 258
rect 1787 250 1791 252
rect 1787 244 1791 246
rect 1787 238 1791 240
rect 1787 232 1791 234
rect 1787 226 1791 228
rect 1787 220 1791 222
rect 1787 214 1791 216
rect 1787 208 1791 210
rect 1787 202 1791 204
rect 1787 196 1791 198
rect 1787 190 1791 192
rect 1787 184 1791 186
rect 1787 178 1791 180
rect 1787 172 1791 174
rect 1787 166 1791 168
rect 1787 160 1791 162
rect 1787 154 1791 156
rect 1787 148 1791 150
rect 2261 508 2265 510
rect 2261 502 2265 504
rect 2261 496 2265 498
rect 2261 490 2265 492
rect 2261 484 2265 486
rect 2261 478 2265 480
rect 2261 472 2265 474
rect 2261 466 2265 468
rect 2261 460 2265 462
rect 2261 454 2265 456
rect 2261 448 2265 450
rect 2261 442 2265 444
rect 2261 436 2265 438
rect 2261 430 2265 432
rect 2261 424 2265 426
rect 2261 418 2265 420
rect 2261 412 2265 414
rect 2261 406 2265 408
rect 2261 400 2265 402
rect 2261 394 2265 396
rect 2261 388 2265 390
rect 2261 382 2265 384
rect 2261 376 2265 378
rect 2261 370 2265 372
rect 2261 364 2265 366
rect 2261 358 2265 360
rect 2261 352 2265 354
rect 2261 346 2265 348
rect 2261 340 2265 342
rect 2261 334 2265 336
rect 2261 328 2265 330
rect 2261 322 2265 324
rect 2261 316 2265 318
rect 2261 310 2265 312
rect 2261 304 2265 306
rect 2261 298 2265 300
rect 2261 292 2265 294
rect 2261 286 2265 288
rect 2261 280 2265 282
rect 2261 274 2265 276
rect 2261 268 2265 270
rect 2261 262 2265 264
rect 2261 256 2265 258
rect 2261 250 2265 252
rect 2261 244 2265 246
rect 2261 238 2265 240
rect 2261 232 2265 234
rect 2261 226 2265 228
rect 2261 220 2265 222
rect 2261 214 2265 216
rect 2261 208 2265 210
rect 2261 202 2265 204
rect 2261 196 2265 198
rect 2261 190 2265 192
rect 2261 184 2265 186
rect 2261 178 2265 180
rect 2261 172 2265 174
rect 2261 166 2265 168
rect 2261 160 2265 162
rect 2261 154 2265 156
rect 2261 148 2265 150
rect 2735 508 2739 510
rect 2735 502 2739 504
rect 2735 496 2739 498
rect 2735 490 2739 492
rect 2735 484 2739 486
rect 2735 478 2739 480
rect 2735 472 2739 474
rect 2735 466 2739 468
rect 2735 460 2739 462
rect 2735 454 2739 456
rect 2735 448 2739 450
rect 2735 442 2739 444
rect 2735 436 2739 438
rect 2735 430 2739 432
rect 2735 424 2739 426
rect 2735 418 2739 420
rect 2735 412 2739 414
rect 2735 406 2739 408
rect 2735 400 2739 402
rect 2735 394 2739 396
rect 2735 388 2739 390
rect 2735 382 2739 384
rect 2735 376 2739 378
rect 2735 370 2739 372
rect 2735 364 2739 366
rect 2735 358 2739 360
rect 2735 352 2739 354
rect 2735 346 2739 348
rect 2735 340 2739 342
rect 2735 334 2739 336
rect 2735 328 2739 330
rect 2735 322 2739 324
rect 2735 316 2739 318
rect 2735 310 2739 312
rect 2735 304 2739 306
rect 2735 298 2739 300
rect 2735 292 2739 294
rect 2735 286 2739 288
rect 2735 280 2739 282
rect 2735 274 2739 276
rect 2735 268 2739 270
rect 2735 262 2739 264
rect 2735 256 2739 258
rect 2735 250 2739 252
rect 2735 244 2739 246
rect 2735 238 2739 240
rect 2735 232 2739 234
rect 2735 226 2739 228
rect 2735 220 2739 222
rect 2735 214 2739 216
rect 2735 208 2739 210
rect 2735 202 2739 204
rect 2735 196 2739 198
rect 2735 190 2739 192
rect 2735 184 2739 186
rect 2735 178 2739 180
rect 2735 172 2739 174
rect 2735 166 2739 168
rect 2735 160 2739 162
rect 2735 154 2739 156
rect 2735 148 2739 150
rect 3209 508 3213 510
rect 3209 502 3213 504
rect 3209 496 3213 498
rect 3209 490 3213 492
rect 3209 484 3213 486
rect 3209 478 3213 480
rect 3209 472 3213 474
rect 3209 466 3213 468
rect 3209 460 3213 462
rect 3209 454 3213 456
rect 3209 448 3213 450
rect 3209 442 3213 444
rect 3209 436 3213 438
rect 3209 430 3213 432
rect 3209 424 3213 426
rect 3209 418 3213 420
rect 3209 412 3213 414
rect 3209 406 3213 408
rect 3209 400 3213 402
rect 3209 394 3213 396
rect 3209 388 3213 390
rect 3209 382 3213 384
rect 3209 376 3213 378
rect 3209 370 3213 372
rect 3209 364 3213 366
rect 3209 358 3213 360
rect 3209 352 3213 354
rect 3209 346 3213 348
rect 3209 340 3213 342
rect 3209 334 3213 336
rect 3209 328 3213 330
rect 3209 322 3213 324
rect 3209 316 3213 318
rect 3209 310 3213 312
rect 3209 304 3213 306
rect 3209 298 3213 300
rect 3209 292 3213 294
rect 3209 286 3213 288
rect 3209 280 3213 282
rect 3209 274 3213 276
rect 3209 268 3213 270
rect 3209 262 3213 264
rect 3209 256 3213 258
rect 3209 250 3213 252
rect 3209 244 3213 246
rect 3209 238 3213 240
rect 3209 232 3213 234
rect 3209 226 3213 228
rect 3209 220 3213 222
rect 3209 214 3213 216
rect 3209 208 3213 210
rect 3209 202 3213 204
rect 3209 196 3213 198
rect 3209 190 3213 192
rect 3209 184 3213 186
rect 3209 178 3213 180
rect 3209 172 3213 174
rect 3209 166 3213 168
rect 3209 160 3213 162
rect 3209 154 3213 156
rect 3209 148 3213 150
rect 3683 508 3687 510
rect 3683 502 3687 504
rect 3683 496 3687 498
rect 3683 490 3687 492
rect 3683 484 3687 486
rect 3683 478 3687 480
rect 3683 472 3687 474
rect 3683 466 3687 468
rect 3683 460 3687 462
rect 3683 454 3687 456
rect 3683 448 3687 450
rect 3683 442 3687 444
rect 3683 436 3687 438
rect 3683 430 3687 432
rect 3683 424 3687 426
rect 3683 418 3687 420
rect 3683 412 3687 414
rect 3683 406 3687 408
rect 3683 400 3687 402
rect 3683 394 3687 396
rect 3683 388 3687 390
rect 3683 382 3687 384
rect 3683 376 3687 378
rect 3683 370 3687 372
rect 3683 364 3687 366
rect 3683 358 3687 360
rect 3683 352 3687 354
rect 3683 346 3687 348
rect 3683 340 3687 342
rect 3683 334 3687 336
rect 3683 328 3687 330
rect 3683 322 3687 324
rect 3683 316 3687 318
rect 3683 310 3687 312
rect 3683 304 3687 306
rect 3683 298 3687 300
rect 3683 292 3687 294
rect 3683 286 3687 288
rect 3683 280 3687 282
rect 3683 274 3687 276
rect 3683 268 3687 270
rect 3683 262 3687 264
rect 3683 256 3687 258
rect 3683 250 3687 252
rect 3683 244 3687 246
rect 3683 238 3687 240
rect 3683 232 3687 234
rect 3683 226 3687 228
rect 3683 220 3687 222
rect 3683 214 3687 216
rect 3683 208 3687 210
rect 3683 202 3687 204
rect 3683 196 3687 198
rect 3683 190 3687 192
rect 3683 184 3687 186
rect 3683 178 3687 180
rect 3683 172 3687 174
rect 3683 166 3687 168
rect 3683 160 3687 162
rect 3683 154 3687 156
rect 3683 148 3687 150
rect 4157 508 4161 510
rect 4157 502 4161 504
rect 4157 496 4161 498
rect 4157 490 4161 492
rect 4157 484 4161 486
rect 4157 478 4161 480
rect 4157 472 4161 474
rect 4157 466 4161 468
rect 4157 460 4161 462
rect 4157 454 4161 456
rect 4157 448 4161 450
rect 4157 442 4161 444
rect 4157 436 4161 438
rect 4157 430 4161 432
rect 4157 424 4161 426
rect 4157 418 4161 420
rect 4157 412 4161 414
rect 4157 406 4161 408
rect 4157 400 4161 402
rect 4157 394 4161 396
rect 4157 388 4161 390
rect 4157 382 4161 384
rect 4157 376 4161 378
rect 4157 370 4161 372
rect 4157 364 4161 366
rect 4157 358 4161 360
rect 4157 352 4161 354
rect 4157 346 4161 348
rect 4157 340 4161 342
rect 4157 334 4161 336
rect 4157 328 4161 330
rect 4157 322 4161 324
rect 4157 316 4161 318
rect 4157 310 4161 312
rect 4157 304 4161 306
rect 4157 298 4161 300
rect 4157 292 4161 294
rect 4157 286 4161 288
rect 4157 280 4161 282
rect 4157 274 4161 276
rect 4157 268 4161 270
rect 4157 262 4161 264
rect 4157 256 4161 258
rect 4157 250 4161 252
rect 4157 244 4161 246
rect 4157 238 4161 240
rect 4157 232 4161 234
rect 4157 226 4161 228
rect 4157 220 4161 222
rect 4157 214 4161 216
rect 4157 208 4161 210
rect 4157 202 4161 204
rect 4157 196 4161 198
rect 4157 190 4161 192
rect 4157 184 4161 186
rect 4157 178 4161 180
rect 4157 172 4161 174
rect 4157 166 4161 168
rect 4157 160 4161 162
rect 4157 154 4161 156
rect 4157 148 4161 150
rect 4631 508 4635 510
rect 4631 502 4635 504
rect 4631 496 4635 498
rect 4631 490 4635 492
rect 4643 499 4684 500
rect 4643 490 4654 499
rect 4668 490 4669 499
rect 4683 490 4684 499
rect 4643 489 4684 490
rect 4631 484 4635 486
rect 4631 478 4635 480
rect 4631 472 4635 474
rect 4631 466 4635 468
rect 4631 460 4635 462
rect 4631 454 4635 456
rect 4631 448 4635 450
rect 4631 442 4635 444
rect 4631 436 4635 438
rect 4631 430 4635 432
rect 4631 424 4635 426
rect 4631 418 4635 420
rect 4631 412 4635 414
rect 4631 406 4635 408
rect 4631 400 4635 402
rect 4631 394 4635 396
rect 4631 388 4635 390
rect 4631 382 4635 384
rect 4631 376 4635 378
rect 4631 370 4635 372
rect 4631 364 4635 366
rect 4631 358 4635 360
rect 4631 352 4635 354
rect 4631 346 4635 348
rect 4631 340 4635 342
rect 4631 334 4635 336
rect 4631 328 4635 330
rect 4631 322 4635 324
rect 4631 316 4635 318
rect 4631 310 4635 312
rect 4631 304 4635 306
rect 4631 298 4635 300
rect 4631 292 4635 294
rect 4631 286 4635 288
rect 4631 280 4635 282
rect 4631 274 4635 276
rect 4631 268 4635 270
rect 4631 262 4635 264
rect 4631 256 4635 258
rect 4631 250 4635 252
rect 4631 244 4635 246
rect 4631 238 4635 240
rect 4631 232 4635 234
rect 4631 226 4635 228
rect 4631 220 4635 222
rect 4631 214 4635 216
rect 4631 208 4635 210
rect 4631 202 4635 204
rect 4673 226 4683 227
rect 4673 212 4674 226
rect 4673 203 4683 212
rect 4631 196 4635 198
rect 4631 190 4635 192
rect 4631 184 4635 186
rect 4653 196 4823 203
rect 4653 190 4813 196
rect 4631 178 4635 180
rect 4631 172 4635 174
rect 4631 166 4635 168
rect 4631 160 4635 162
rect 4653 176 4669 190
rect 4657 172 4659 176
rect 4663 172 4665 176
rect 4653 170 4669 172
rect 4657 166 4659 170
rect 4663 166 4665 170
rect 4647 156 4651 160
rect 4671 156 4675 160
rect 4687 180 4691 182
rect 4687 174 4691 176
rect 4687 168 4691 170
rect 4687 162 4691 164
rect 4687 156 4691 158
rect 4709 176 4725 190
rect 4753 188 4763 190
rect 4713 172 4715 176
rect 4719 172 4721 176
rect 4709 170 4725 172
rect 4713 166 4715 170
rect 4719 166 4721 170
rect 4703 156 4707 160
rect 4727 156 4731 160
rect 4743 180 4747 182
rect 4743 174 4747 176
rect 4743 168 4747 170
rect 4743 162 4747 164
rect 4743 156 4747 158
rect 4631 154 4635 156
rect 4631 148 4635 150
rect 4687 148 4691 152
rect 4757 184 4759 188
rect 4779 188 4789 190
rect 4753 182 4763 184
rect 4757 178 4759 182
rect 4753 176 4763 178
rect 4757 172 4759 176
rect 4753 170 4763 172
rect 4757 166 4759 170
rect 4753 164 4763 166
rect 4757 160 4759 164
rect 4753 158 4763 160
rect 4757 154 4759 158
rect 4769 180 4773 182
rect 4769 174 4773 176
rect 4769 168 4773 170
rect 4769 162 4773 164
rect 4769 156 4773 158
rect 4743 148 4747 152
rect 4783 184 4785 188
rect 4779 182 4789 184
rect 4783 178 4785 182
rect 4779 176 4789 178
rect 4783 172 4785 176
rect 4779 170 4789 172
rect 4783 166 4785 170
rect 4779 164 4789 166
rect 4783 160 4785 164
rect 4779 158 4789 160
rect 4783 154 4785 158
rect 4795 180 4799 182
rect 4812 182 4813 190
rect 4822 182 4823 196
rect 4971 196 4987 253
rect 4971 187 4972 196
rect 4986 187 4987 196
rect 4971 186 4987 187
rect 4812 181 4823 182
rect 4795 174 4799 176
rect 4795 168 4799 170
rect 4795 162 4799 164
rect 4795 156 4799 158
rect 4769 148 4773 152
rect 4795 148 4799 152
rect 3 144 5 148
rect 9 144 11 148
rect 15 144 17 148
rect 21 144 23 148
rect 27 144 29 148
rect 33 144 35 148
rect 39 144 41 148
rect 45 144 47 148
rect 51 144 53 148
rect 57 144 59 148
rect 63 144 65 148
rect 69 144 71 148
rect 75 144 77 148
rect 81 144 83 148
rect 87 144 89 148
rect 93 144 95 148
rect 99 144 101 148
rect 105 144 107 148
rect 111 144 113 148
rect 117 144 119 148
rect 123 144 125 148
rect 129 144 131 148
rect 135 144 137 148
rect 141 144 143 148
rect 147 144 149 148
rect 153 144 155 148
rect 159 144 161 148
rect 165 144 167 148
rect 171 144 173 148
rect 177 144 179 148
rect 183 144 185 148
rect 189 144 191 148
rect 195 144 197 148
rect 201 144 203 148
rect 207 144 209 148
rect 213 144 215 148
rect 219 144 221 148
rect 225 144 227 148
rect 231 144 233 148
rect 237 144 239 148
rect 243 144 245 148
rect 249 144 251 148
rect 255 144 257 148
rect 261 144 263 148
rect 267 144 269 148
rect 273 144 275 148
rect 279 144 281 148
rect 285 144 287 148
rect 291 144 293 148
rect 297 144 299 148
rect 303 144 305 148
rect 309 144 311 148
rect 315 144 317 148
rect 321 144 323 148
rect 327 144 329 148
rect 333 144 335 148
rect 339 144 341 148
rect 345 144 347 148
rect 351 144 353 148
rect 357 144 359 148
rect 363 144 365 148
rect 369 144 371 148
rect 375 144 377 148
rect 381 144 383 148
rect 387 144 389 148
rect 393 144 395 148
rect 399 144 401 148
rect 405 144 407 148
rect 411 144 413 148
rect 417 144 419 148
rect 423 144 425 148
rect 429 144 431 148
rect 435 144 437 148
rect 441 144 443 148
rect 447 144 449 148
rect 453 144 455 148
rect 459 144 461 148
rect 465 144 467 148
rect 471 144 473 148
rect 477 144 479 148
rect 483 144 485 148
rect 489 144 491 148
rect 495 144 497 148
rect 501 144 503 148
rect 507 144 509 148
rect 513 144 515 148
rect 519 144 521 148
rect 525 144 527 148
rect 531 144 533 148
rect 537 144 539 148
rect 543 144 545 148
rect 549 144 551 148
rect 555 144 557 148
rect 561 144 563 148
rect 567 144 569 148
rect 573 144 575 148
rect 579 144 581 148
rect 585 144 587 148
rect 621 144 623 148
rect 627 144 629 148
rect 633 144 635 148
rect 639 144 641 148
rect 645 144 647 148
rect 651 144 653 148
rect 657 144 659 148
rect 663 144 665 148
rect 669 144 671 148
rect 675 144 677 148
rect 681 144 683 148
rect 687 144 689 148
rect 693 144 695 148
rect 699 144 701 148
rect 705 144 707 148
rect 711 144 713 148
rect 717 144 719 148
rect 723 144 725 148
rect 729 144 731 148
rect 735 144 737 148
rect 741 144 743 148
rect 747 144 749 148
rect 753 144 755 148
rect 759 144 761 148
rect 765 144 767 148
rect 771 144 773 148
rect 777 144 779 148
rect 783 144 785 148
rect 789 144 791 148
rect 795 144 797 148
rect 801 144 803 148
rect 807 144 809 148
rect 813 144 815 148
rect 819 144 821 148
rect 825 144 827 148
rect 831 144 833 148
rect 837 144 839 148
rect 843 144 845 148
rect 849 144 851 148
rect 855 144 857 148
rect 861 144 863 148
rect 867 144 869 148
rect 873 144 875 148
rect 879 144 881 148
rect 885 144 887 148
rect 891 144 893 148
rect 897 144 899 148
rect 903 144 905 148
rect 909 144 911 148
rect 915 144 917 148
rect 921 144 923 148
rect 927 144 929 148
rect 933 144 935 148
rect 939 144 941 148
rect 945 144 947 148
rect 951 144 953 148
rect 957 144 959 148
rect 963 144 965 148
rect 969 144 971 148
rect 975 144 977 148
rect 981 144 983 148
rect 987 144 989 148
rect 993 144 995 148
rect 999 144 1001 148
rect 1005 144 1007 148
rect 1011 144 1013 148
rect 1017 144 1019 148
rect 1023 144 1025 148
rect 1029 144 1031 148
rect 1035 144 1037 148
rect 1041 144 1043 148
rect 1047 144 1049 148
rect 1053 144 1055 148
rect 1059 144 1061 148
rect 1095 144 1097 148
rect 1101 144 1103 148
rect 1107 144 1109 148
rect 1113 144 1115 148
rect 1119 144 1121 148
rect 1125 144 1127 148
rect 1131 144 1133 148
rect 1137 144 1139 148
rect 1143 144 1145 148
rect 1149 144 1151 148
rect 1155 144 1157 148
rect 1161 144 1163 148
rect 1167 144 1169 148
rect 1173 144 1175 148
rect 1179 144 1181 148
rect 1185 144 1187 148
rect 1191 144 1193 148
rect 1197 144 1199 148
rect 1203 144 1205 148
rect 1209 144 1211 148
rect 1215 144 1217 148
rect 1221 144 1223 148
rect 1227 144 1229 148
rect 1233 144 1235 148
rect 1239 144 1241 148
rect 1245 144 1247 148
rect 1251 144 1253 148
rect 1257 144 1259 148
rect 1263 144 1265 148
rect 1269 144 1271 148
rect 1275 144 1277 148
rect 1281 144 1283 148
rect 1287 144 1289 148
rect 1293 144 1295 148
rect 1299 144 1301 148
rect 1305 144 1307 148
rect 1311 144 1313 148
rect 1317 144 1319 148
rect 1323 144 1325 148
rect 1329 144 1331 148
rect 1335 144 1337 148
rect 1341 144 1343 148
rect 1347 144 1349 148
rect 1353 144 1355 148
rect 1359 144 1361 148
rect 1365 144 1367 148
rect 1371 144 1373 148
rect 1377 144 1379 148
rect 1383 144 1385 148
rect 1389 144 1391 148
rect 1395 144 1397 148
rect 1401 144 1403 148
rect 1407 144 1409 148
rect 1413 144 1415 148
rect 1419 144 1421 148
rect 1425 144 1427 148
rect 1431 144 1433 148
rect 1437 144 1439 148
rect 1443 144 1445 148
rect 1449 144 1451 148
rect 1455 144 1457 148
rect 1461 144 1463 148
rect 1467 144 1469 148
rect 1473 144 1475 148
rect 1479 144 1481 148
rect 1485 144 1487 148
rect 1491 144 1493 148
rect 1497 144 1499 148
rect 1503 144 1505 148
rect 1509 144 1511 148
rect 1515 144 1517 148
rect 1521 144 1523 148
rect 1527 144 1529 148
rect 1533 144 1535 148
rect 1569 144 1571 148
rect 1575 144 1577 148
rect 1581 144 1583 148
rect 1587 144 1589 148
rect 1593 144 1595 148
rect 1599 144 1601 148
rect 1605 144 1607 148
rect 1611 144 1613 148
rect 1617 144 1619 148
rect 1623 144 1625 148
rect 1629 144 1631 148
rect 1635 144 1637 148
rect 1641 144 1643 148
rect 1647 144 1649 148
rect 1653 144 1655 148
rect 1659 144 1661 148
rect 1665 144 1667 148
rect 1671 144 1673 148
rect 1677 144 1679 148
rect 1683 144 1685 148
rect 1689 144 1691 148
rect 1695 144 1697 148
rect 1701 144 1703 148
rect 1707 144 1709 148
rect 1713 144 1715 148
rect 1719 144 1721 148
rect 1725 144 1727 148
rect 1731 144 1733 148
rect 1737 144 1739 148
rect 1743 144 1745 148
rect 1749 144 1751 148
rect 1755 144 1757 148
rect 1761 144 1763 148
rect 1767 144 1769 148
rect 1773 144 1775 148
rect 1779 144 1781 148
rect 1785 144 1787 148
rect 1791 144 1793 148
rect 1797 144 1799 148
rect 1803 144 1805 148
rect 1809 144 1811 148
rect 1815 144 1817 148
rect 1821 144 1823 148
rect 1827 144 1829 148
rect 1833 144 1835 148
rect 1839 144 1841 148
rect 1845 144 1847 148
rect 1851 144 1853 148
rect 1857 144 1859 148
rect 1863 144 1865 148
rect 1869 144 1871 148
rect 1875 144 1877 148
rect 1881 144 1883 148
rect 1887 144 1889 148
rect 1893 144 1895 148
rect 1899 144 1901 148
rect 1905 144 1907 148
rect 1911 144 1913 148
rect 1917 144 1919 148
rect 1923 144 1925 148
rect 1929 144 1931 148
rect 1935 144 1937 148
rect 1941 144 1943 148
rect 1947 144 1949 148
rect 1953 144 1955 148
rect 1959 144 1961 148
rect 1965 144 1967 148
rect 1971 144 1973 148
rect 1977 144 1979 148
rect 1983 144 1985 148
rect 1989 144 1991 148
rect 1995 144 1997 148
rect 2001 144 2003 148
rect 2007 144 2009 148
rect 2043 144 2045 148
rect 2049 144 2051 148
rect 2055 144 2057 148
rect 2061 144 2063 148
rect 2067 144 2069 148
rect 2073 144 2075 148
rect 2079 144 2081 148
rect 2085 144 2087 148
rect 2091 144 2093 148
rect 2097 144 2099 148
rect 2103 144 2105 148
rect 2109 144 2111 148
rect 2115 144 2117 148
rect 2121 144 2123 148
rect 2127 144 2129 148
rect 2133 144 2135 148
rect 2139 144 2141 148
rect 2145 144 2147 148
rect 2151 144 2153 148
rect 2157 144 2159 148
rect 2163 144 2165 148
rect 2169 144 2171 148
rect 2175 144 2177 148
rect 2181 144 2183 148
rect 2187 144 2189 148
rect 2193 144 2195 148
rect 2199 144 2201 148
rect 2205 144 2207 148
rect 2211 144 2213 148
rect 2217 144 2219 148
rect 2223 144 2225 148
rect 2229 144 2231 148
rect 2235 144 2237 148
rect 2241 144 2243 148
rect 2247 144 2249 148
rect 2253 144 2255 148
rect 2259 144 2261 148
rect 2265 144 2267 148
rect 2271 144 2273 148
rect 2277 144 2279 148
rect 2283 144 2285 148
rect 2289 144 2291 148
rect 2295 144 2297 148
rect 2301 144 2303 148
rect 2307 144 2309 148
rect 2313 144 2315 148
rect 2319 144 2321 148
rect 2325 144 2327 148
rect 2331 144 2333 148
rect 2337 144 2339 148
rect 2343 144 2345 148
rect 2349 144 2351 148
rect 2355 144 2357 148
rect 2361 144 2363 148
rect 2367 144 2369 148
rect 2373 144 2375 148
rect 2379 144 2381 148
rect 2385 144 2387 148
rect 2391 144 2393 148
rect 2397 144 2399 148
rect 2403 144 2405 148
rect 2409 144 2411 148
rect 2415 144 2417 148
rect 2421 144 2423 148
rect 2427 144 2429 148
rect 2433 144 2435 148
rect 2439 144 2441 148
rect 2445 144 2447 148
rect 2451 144 2453 148
rect 2457 144 2459 148
rect 2463 144 2465 148
rect 2469 144 2471 148
rect 2475 144 2477 148
rect 2481 144 2483 148
rect 2517 144 2519 148
rect 2523 144 2525 148
rect 2529 144 2531 148
rect 2535 144 2537 148
rect 2541 144 2543 148
rect 2547 144 2549 148
rect 2553 144 2555 148
rect 2559 144 2561 148
rect 2565 144 2567 148
rect 2571 144 2573 148
rect 2577 144 2579 148
rect 2583 144 2585 148
rect 2589 144 2591 148
rect 2595 144 2597 148
rect 2601 144 2603 148
rect 2607 144 2609 148
rect 2613 144 2615 148
rect 2619 144 2621 148
rect 2625 144 2627 148
rect 2631 144 2633 148
rect 2637 144 2639 148
rect 2643 144 2645 148
rect 2649 144 2651 148
rect 2655 144 2657 148
rect 2661 144 2663 148
rect 2667 144 2669 148
rect 2673 144 2675 148
rect 2679 144 2681 148
rect 2685 144 2687 148
rect 2691 144 2693 148
rect 2697 144 2699 148
rect 2703 144 2705 148
rect 2709 144 2711 148
rect 2715 144 2717 148
rect 2721 144 2723 148
rect 2727 144 2729 148
rect 2733 144 2735 148
rect 2739 144 2741 148
rect 2745 144 2747 148
rect 2751 144 2753 148
rect 2757 144 2759 148
rect 2763 144 2765 148
rect 2769 144 2771 148
rect 2775 144 2777 148
rect 2781 144 2783 148
rect 2787 144 2789 148
rect 2793 144 2795 148
rect 2799 144 2801 148
rect 2805 144 2807 148
rect 2811 144 2813 148
rect 2817 144 2819 148
rect 2823 144 2825 148
rect 2829 144 2831 148
rect 2835 144 2837 148
rect 2841 144 2843 148
rect 2847 144 2849 148
rect 2853 144 2855 148
rect 2859 144 2861 148
rect 2865 144 2867 148
rect 2871 144 2873 148
rect 2877 144 2879 148
rect 2883 144 2885 148
rect 2889 144 2891 148
rect 2895 144 2897 148
rect 2901 144 2903 148
rect 2907 144 2909 148
rect 2913 144 2915 148
rect 2919 144 2921 148
rect 2925 144 2927 148
rect 2931 144 2933 148
rect 2937 144 2939 148
rect 2943 144 2945 148
rect 2949 144 2951 148
rect 2955 144 2957 148
rect 2991 144 2993 148
rect 2997 144 2999 148
rect 3003 144 3005 148
rect 3009 144 3011 148
rect 3015 144 3017 148
rect 3021 144 3023 148
rect 3027 144 3029 148
rect 3033 144 3035 148
rect 3039 144 3041 148
rect 3045 144 3047 148
rect 3051 144 3053 148
rect 3057 144 3059 148
rect 3063 144 3065 148
rect 3069 144 3071 148
rect 3075 144 3077 148
rect 3081 144 3083 148
rect 3087 144 3089 148
rect 3093 144 3095 148
rect 3099 144 3101 148
rect 3105 144 3107 148
rect 3111 144 3113 148
rect 3117 144 3119 148
rect 3123 144 3125 148
rect 3129 144 3131 148
rect 3135 144 3137 148
rect 3141 144 3143 148
rect 3147 144 3149 148
rect 3153 144 3155 148
rect 3159 144 3161 148
rect 3165 144 3167 148
rect 3171 144 3173 148
rect 3177 144 3179 148
rect 3183 144 3185 148
rect 3189 144 3191 148
rect 3195 144 3197 148
rect 3201 144 3203 148
rect 3207 144 3209 148
rect 3213 144 3215 148
rect 3219 144 3221 148
rect 3225 144 3227 148
rect 3231 144 3233 148
rect 3237 144 3239 148
rect 3243 144 3245 148
rect 3249 144 3251 148
rect 3255 144 3257 148
rect 3261 144 3263 148
rect 3267 144 3269 148
rect 3273 144 3275 148
rect 3279 144 3281 148
rect 3285 144 3287 148
rect 3291 144 3293 148
rect 3297 144 3299 148
rect 3303 144 3305 148
rect 3309 144 3311 148
rect 3315 144 3317 148
rect 3321 144 3323 148
rect 3327 144 3329 148
rect 3333 144 3335 148
rect 3339 144 3341 148
rect 3345 144 3347 148
rect 3351 144 3353 148
rect 3357 144 3359 148
rect 3363 144 3365 148
rect 3369 144 3371 148
rect 3375 144 3377 148
rect 3381 144 3383 148
rect 3387 144 3389 148
rect 3393 144 3395 148
rect 3399 144 3401 148
rect 3405 144 3407 148
rect 3411 144 3413 148
rect 3417 144 3419 148
rect 3423 144 3425 148
rect 3429 144 3431 148
rect 3465 144 3467 148
rect 3471 144 3473 148
rect 3477 144 3479 148
rect 3483 144 3485 148
rect 3489 144 3491 148
rect 3495 144 3497 148
rect 3501 144 3503 148
rect 3507 144 3509 148
rect 3513 144 3515 148
rect 3519 144 3521 148
rect 3525 144 3527 148
rect 3531 144 3533 148
rect 3537 144 3539 148
rect 3543 144 3545 148
rect 3549 144 3551 148
rect 3555 144 3557 148
rect 3561 144 3563 148
rect 3567 144 3569 148
rect 3573 144 3575 148
rect 3579 144 3581 148
rect 3585 144 3587 148
rect 3591 144 3593 148
rect 3597 144 3599 148
rect 3603 144 3605 148
rect 3609 144 3611 148
rect 3615 144 3617 148
rect 3621 144 3623 148
rect 3627 144 3629 148
rect 3633 144 3635 148
rect 3639 144 3641 148
rect 3645 144 3647 148
rect 3651 144 3653 148
rect 3657 144 3659 148
rect 3663 144 3665 148
rect 3669 144 3671 148
rect 3675 144 3677 148
rect 3681 144 3683 148
rect 3687 144 3689 148
rect 3693 144 3695 148
rect 3699 144 3701 148
rect 3705 144 3707 148
rect 3711 144 3713 148
rect 3717 144 3719 148
rect 3723 144 3725 148
rect 3729 144 3731 148
rect 3735 144 3737 148
rect 3741 144 3743 148
rect 3747 144 3749 148
rect 3753 144 3755 148
rect 3759 144 3761 148
rect 3765 144 3767 148
rect 3771 144 3773 148
rect 3777 144 3779 148
rect 3783 144 3785 148
rect 3789 144 3791 148
rect 3795 144 3797 148
rect 3801 144 3803 148
rect 3807 144 3809 148
rect 3813 144 3815 148
rect 3819 144 3821 148
rect 3825 144 3827 148
rect 3831 144 3833 148
rect 3837 144 3839 148
rect 3843 144 3845 148
rect 3849 144 3851 148
rect 3855 144 3857 148
rect 3861 144 3863 148
rect 3867 144 3869 148
rect 3873 144 3875 148
rect 3879 144 3881 148
rect 3885 144 3887 148
rect 3891 144 3893 148
rect 3897 144 3899 148
rect 3903 144 3905 148
rect 3939 144 3941 148
rect 3945 144 3947 148
rect 3951 144 3953 148
rect 3957 144 3959 148
rect 3963 144 3965 148
rect 3969 144 3971 148
rect 3975 144 3977 148
rect 3981 144 3983 148
rect 3987 144 3989 148
rect 3993 144 3995 148
rect 3999 144 4001 148
rect 4005 144 4007 148
rect 4011 144 4013 148
rect 4017 144 4019 148
rect 4023 144 4025 148
rect 4029 144 4031 148
rect 4035 144 4037 148
rect 4041 144 4043 148
rect 4047 144 4049 148
rect 4053 144 4055 148
rect 4059 144 4061 148
rect 4065 144 4067 148
rect 4071 144 4073 148
rect 4077 144 4079 148
rect 4083 144 4085 148
rect 4089 144 4091 148
rect 4095 144 4097 148
rect 4101 144 4103 148
rect 4107 144 4109 148
rect 4113 144 4115 148
rect 4119 144 4121 148
rect 4125 144 4127 148
rect 4131 144 4133 148
rect 4137 144 4139 148
rect 4143 144 4145 148
rect 4149 144 4151 148
rect 4155 144 4157 148
rect 4161 144 4163 148
rect 4167 144 4169 148
rect 4173 144 4175 148
rect 4179 144 4181 148
rect 4185 144 4187 148
rect 4191 144 4193 148
rect 4197 144 4199 148
rect 4203 144 4205 148
rect 4209 144 4211 148
rect 4215 144 4217 148
rect 4221 144 4223 148
rect 4227 144 4229 148
rect 4233 144 4235 148
rect 4239 144 4241 148
rect 4245 144 4247 148
rect 4251 144 4253 148
rect 4257 144 4259 148
rect 4263 144 4265 148
rect 4269 144 4271 148
rect 4275 144 4277 148
rect 4281 144 4283 148
rect 4287 144 4289 148
rect 4293 144 4295 148
rect 4299 144 4301 148
rect 4305 144 4307 148
rect 4311 144 4313 148
rect 4317 144 4319 148
rect 4323 144 4325 148
rect 4329 144 4331 148
rect 4335 144 4337 148
rect 4341 144 4343 148
rect 4347 144 4349 148
rect 4353 144 4355 148
rect 4359 144 4361 148
rect 4365 144 4367 148
rect 4371 144 4373 148
rect 4377 144 4379 148
rect 4413 144 4415 148
rect 4419 144 4421 148
rect 4425 144 4427 148
rect 4431 144 4433 148
rect 4437 144 4439 148
rect 4443 144 4445 148
rect 4449 144 4451 148
rect 4455 144 4457 148
rect 4461 144 4463 148
rect 4467 144 4469 148
rect 4473 144 4475 148
rect 4479 144 4481 148
rect 4485 144 4487 148
rect 4491 144 4493 148
rect 4497 144 4499 148
rect 4503 144 4505 148
rect 4509 144 4511 148
rect 4515 144 4517 148
rect 4521 144 4523 148
rect 4527 144 4529 148
rect 4533 144 4535 148
rect 4539 144 4541 148
rect 4545 144 4547 148
rect 4551 144 4553 148
rect 4557 144 4559 148
rect 4563 144 4565 148
rect 4569 144 4571 148
rect 4575 144 4577 148
rect 4581 144 4583 148
rect 4587 144 4589 148
rect 4593 144 4595 148
rect 4599 144 4601 148
rect 4605 144 4607 148
rect 4611 144 4613 148
rect 4617 144 4619 148
rect 4623 144 4625 148
rect 4629 144 4631 148
rect 4635 144 4637 148
rect 4641 144 4643 148
rect 4647 144 4649 148
rect 4653 144 4655 148
rect 4659 144 4661 148
rect 4665 144 4667 148
rect 4671 144 4673 148
rect 4677 144 4679 148
rect 4683 144 4685 148
rect 4689 144 4691 148
rect 4695 144 4697 148
rect 4701 144 4703 148
rect 4707 144 4709 148
rect 4713 144 4715 148
rect 4719 144 4721 148
rect 4725 144 4727 148
rect 4731 144 4733 148
rect 4737 144 4739 148
rect 4743 144 4745 148
rect 4749 144 4751 148
rect 4755 144 4757 148
rect 4761 144 4763 148
rect 4767 144 4769 148
rect 4773 144 4775 148
rect 4779 144 4781 148
rect 4785 144 4787 148
rect 4791 144 4793 148
rect 4797 144 4799 148
rect 4803 144 4805 148
rect 4809 144 4811 148
rect 4815 144 4817 148
rect 4821 144 4823 148
rect 4827 144 4829 148
rect 4833 144 4835 148
rect 4839 144 4841 148
rect 4845 144 4847 148
rect 4851 144 4853 148
rect 4857 144 4859 148
rect 4863 144 4865 148
rect 4869 144 4871 148
rect 4875 144 4877 148
rect 4881 144 4883 148
rect 4887 144 4889 148
rect 4893 144 4895 148
rect 4899 144 4901 148
rect 4905 144 4907 148
rect 4911 144 4913 148
rect 4917 144 4919 148
rect 4923 144 4925 148
rect 4929 144 4931 148
rect 4935 144 4937 148
rect 4941 144 4943 148
rect 4947 144 4949 148
rect 4953 144 4955 148
rect 4959 144 4961 148
rect 4965 144 4967 148
rect 4971 144 4973 148
rect 4977 144 4979 148
rect 4983 144 4985 148
rect 4989 144 4991 148
rect 4995 144 4997 148
rect 495 141 535 144
rect 499 137 501 141
rect 505 137 507 141
rect 511 137 513 141
rect 517 137 519 141
rect 523 137 525 141
rect 529 137 531 141
rect 495 101 535 137
rect 673 141 713 144
rect 677 137 679 141
rect 683 137 685 141
rect 689 137 691 141
rect 695 137 697 141
rect 701 137 703 141
rect 707 137 709 141
rect 549 131 551 135
rect 555 131 557 135
rect 561 131 563 135
rect 567 131 569 135
rect 573 131 575 135
rect 545 129 579 131
rect 543 125 545 129
rect 549 125 551 129
rect 555 125 557 129
rect 561 125 563 129
rect 567 125 569 129
rect 573 125 575 129
rect 539 123 579 125
rect 543 119 545 123
rect 549 119 551 123
rect 555 119 557 123
rect 561 119 563 123
rect 567 119 569 123
rect 573 119 575 123
rect 539 116 579 119
rect 543 112 545 116
rect 549 112 551 116
rect 555 112 557 116
rect 561 112 563 116
rect 567 112 569 116
rect 573 112 575 116
rect 539 111 579 112
rect 543 107 545 111
rect 549 107 551 111
rect 555 107 557 111
rect 561 107 563 111
rect 567 107 569 111
rect 573 107 575 111
rect 633 131 635 135
rect 639 131 641 135
rect 645 131 647 135
rect 651 131 653 135
rect 657 131 659 135
rect 629 129 663 131
rect 633 125 635 129
rect 639 125 641 129
rect 645 125 647 129
rect 651 125 653 129
rect 657 125 659 129
rect 663 125 665 129
rect 629 123 669 125
rect 633 119 635 123
rect 639 119 641 123
rect 645 119 647 123
rect 651 119 653 123
rect 657 119 659 123
rect 663 119 665 123
rect 629 116 669 119
rect 633 112 635 116
rect 639 112 641 116
rect 645 112 647 116
rect 651 112 653 116
rect 657 112 659 116
rect 663 112 665 116
rect 629 111 669 112
rect 633 107 635 111
rect 639 107 641 111
rect 645 107 647 111
rect 651 107 653 111
rect 657 107 659 111
rect 663 107 665 111
rect 499 92 501 101
rect 505 92 507 101
rect 511 92 513 101
rect 517 92 519 101
rect 523 92 525 101
rect 529 92 531 101
rect 673 101 713 137
rect 495 90 535 92
rect 499 86 501 90
rect 505 86 507 90
rect 511 86 513 90
rect 517 86 519 90
rect 523 86 525 90
rect 529 86 531 90
rect 495 84 535 86
rect 499 80 501 84
rect 505 80 507 84
rect 511 80 513 84
rect 517 80 519 84
rect 523 80 525 84
rect 529 80 531 84
rect 495 78 535 80
rect 499 74 501 78
rect 505 74 507 78
rect 511 74 513 78
rect 517 74 519 78
rect 523 74 525 78
rect 529 74 531 78
rect 495 72 535 74
rect 499 63 501 72
rect 505 63 507 72
rect 511 63 513 72
rect 517 63 519 72
rect 523 63 525 72
rect 529 63 531 72
rect 495 62 535 63
rect 539 99 569 100
rect 539 95 540 99
rect 544 95 546 99
rect 550 95 552 99
rect 556 95 558 99
rect 562 95 564 99
rect 568 95 569 99
rect 539 93 569 95
rect 539 89 540 93
rect 544 89 546 93
rect 550 89 552 93
rect 556 89 558 93
rect 562 89 564 93
rect 568 89 569 93
rect 539 86 569 89
rect 539 82 540 86
rect 544 82 546 86
rect 550 82 552 86
rect 556 82 558 86
rect 562 82 564 86
rect 568 82 569 86
rect 539 80 569 82
rect 539 76 540 80
rect 544 76 546 80
rect 550 76 552 80
rect 556 76 558 80
rect 562 76 564 80
rect 568 76 569 80
rect 539 74 569 76
rect 539 70 540 74
rect 544 70 546 74
rect 550 70 552 74
rect 556 70 558 74
rect 562 70 564 74
rect 568 70 569 74
rect 539 68 569 70
rect 539 64 540 68
rect 544 64 546 68
rect 550 64 552 68
rect 556 64 558 68
rect 562 64 564 68
rect 568 64 569 68
rect 539 48 569 64
rect 639 99 669 100
rect 639 95 640 99
rect 644 95 646 99
rect 650 95 652 99
rect 656 95 658 99
rect 662 95 664 99
rect 668 95 669 99
rect 639 93 669 95
rect 639 89 640 93
rect 644 89 646 93
rect 650 89 652 93
rect 656 89 658 93
rect 662 89 664 93
rect 668 89 669 93
rect 639 86 669 89
rect 639 82 640 86
rect 644 82 646 86
rect 650 82 652 86
rect 656 82 658 86
rect 662 82 664 86
rect 668 82 669 86
rect 639 80 669 82
rect 639 76 640 80
rect 644 76 646 80
rect 650 76 652 80
rect 656 76 658 80
rect 662 76 664 80
rect 668 76 669 80
rect 639 74 669 76
rect 639 70 640 74
rect 644 70 646 74
rect 650 70 652 74
rect 656 70 658 74
rect 662 70 664 74
rect 668 70 669 74
rect 639 68 669 70
rect 639 64 640 68
rect 644 64 646 68
rect 650 64 652 68
rect 656 64 658 68
rect 662 64 664 68
rect 668 64 669 68
rect 573 57 592 58
rect 577 53 578 57
rect 582 53 583 57
rect 587 53 588 57
rect 573 52 592 53
rect 539 47 579 48
rect 543 43 545 47
rect 549 43 551 47
rect 555 43 557 47
rect 561 43 563 47
rect 567 43 569 47
rect 573 43 575 47
rect 539 42 579 43
rect 543 38 545 42
rect 549 38 551 42
rect 555 38 557 42
rect 561 38 563 42
rect 567 38 569 42
rect 573 38 575 42
rect 539 36 579 38
rect 543 32 545 36
rect 549 32 551 36
rect 555 32 557 36
rect 561 32 563 36
rect 567 32 569 36
rect 573 32 575 36
rect 539 30 579 32
rect 543 26 545 30
rect 549 26 551 30
rect 555 26 557 30
rect 561 26 563 30
rect 567 26 569 30
rect 573 26 575 30
rect 539 24 579 26
rect 543 20 545 24
rect 549 20 551 24
rect 555 20 557 24
rect 561 20 563 24
rect 567 20 569 24
rect 573 20 575 24
rect 539 18 579 20
rect 543 14 545 18
rect 549 14 551 18
rect 555 14 557 18
rect 561 14 563 18
rect 567 14 569 18
rect 573 14 575 18
rect 539 4 579 14
rect 543 0 545 4
rect 549 0 551 4
rect 555 0 557 4
rect 561 0 563 4
rect 567 0 569 4
rect 573 0 575 4
rect 583 4 592 52
rect 616 57 635 58
rect 620 53 621 57
rect 625 53 626 57
rect 630 53 631 57
rect 616 52 635 53
rect 616 4 625 52
rect 639 48 669 64
rect 629 47 669 48
rect 633 43 635 47
rect 639 43 641 47
rect 645 43 647 47
rect 651 43 653 47
rect 657 43 659 47
rect 663 43 665 47
rect 629 42 669 43
rect 633 38 635 42
rect 639 38 641 42
rect 645 38 647 42
rect 651 38 653 42
rect 657 38 659 42
rect 663 38 665 42
rect 629 36 669 38
rect 633 32 635 36
rect 639 32 641 36
rect 645 32 647 36
rect 651 32 653 36
rect 657 32 659 36
rect 663 32 665 36
rect 629 30 669 32
rect 633 26 635 30
rect 639 26 641 30
rect 645 26 647 30
rect 651 26 653 30
rect 657 26 659 30
rect 663 26 665 30
rect 629 24 669 26
rect 633 20 635 24
rect 639 20 641 24
rect 645 20 647 24
rect 651 20 653 24
rect 657 20 659 24
rect 663 20 665 24
rect 629 18 669 20
rect 633 14 635 18
rect 639 14 641 18
rect 645 14 647 18
rect 651 14 653 18
rect 657 14 659 18
rect 663 14 669 18
rect 629 4 669 14
rect 633 0 635 4
rect 639 0 641 4
rect 645 0 647 4
rect 651 0 653 4
rect 657 0 659 4
rect 663 0 665 4
rect 677 92 679 101
rect 683 92 685 101
rect 689 92 691 101
rect 695 92 697 101
rect 701 92 703 101
rect 707 92 709 101
rect 673 90 713 92
rect 677 86 679 90
rect 683 86 685 90
rect 689 86 691 90
rect 695 86 697 90
rect 701 86 703 90
rect 707 86 709 90
rect 673 84 713 86
rect 677 80 679 84
rect 683 80 685 84
rect 689 80 691 84
rect 695 80 697 84
rect 701 80 703 84
rect 707 80 709 84
rect 673 78 713 80
rect 677 74 679 78
rect 683 74 685 78
rect 689 74 691 78
rect 695 74 697 78
rect 701 74 703 78
rect 707 74 709 78
rect 673 72 713 74
rect 677 63 679 72
rect 683 63 685 72
rect 689 63 691 72
rect 695 63 697 72
rect 701 63 703 72
rect 707 63 709 72
rect 673 12 713 63
rect 677 8 679 12
rect 683 8 685 12
rect 689 8 691 12
rect 695 8 697 12
rect 701 8 703 12
rect 707 8 709 12
rect 673 4 713 8
rect 677 0 679 4
rect 683 0 685 4
rect 689 0 691 4
rect 695 0 697 4
rect 701 0 703 4
rect 707 0 709 4
rect 969 141 1009 144
rect 973 137 975 141
rect 979 137 981 141
rect 985 137 987 141
rect 991 137 993 141
rect 997 137 999 141
rect 1003 137 1005 141
rect 969 101 1009 137
rect 1147 141 1187 144
rect 1151 137 1153 141
rect 1157 137 1159 141
rect 1163 137 1165 141
rect 1169 137 1171 141
rect 1175 137 1177 141
rect 1181 137 1183 141
rect 1023 131 1025 135
rect 1029 131 1031 135
rect 1035 131 1037 135
rect 1041 131 1043 135
rect 1047 131 1049 135
rect 1019 129 1053 131
rect 1017 125 1019 129
rect 1023 125 1025 129
rect 1029 125 1031 129
rect 1035 125 1037 129
rect 1041 125 1043 129
rect 1047 125 1049 129
rect 1013 123 1053 125
rect 1017 119 1019 123
rect 1023 119 1025 123
rect 1029 119 1031 123
rect 1035 119 1037 123
rect 1041 119 1043 123
rect 1047 119 1049 123
rect 1013 116 1053 119
rect 1017 112 1019 116
rect 1023 112 1025 116
rect 1029 112 1031 116
rect 1035 112 1037 116
rect 1041 112 1043 116
rect 1047 112 1049 116
rect 1013 111 1053 112
rect 1017 107 1019 111
rect 1023 107 1025 111
rect 1029 107 1031 111
rect 1035 107 1037 111
rect 1041 107 1043 111
rect 1047 107 1049 111
rect 1107 131 1109 135
rect 1113 131 1115 135
rect 1119 131 1121 135
rect 1125 131 1127 135
rect 1131 131 1133 135
rect 1103 129 1137 131
rect 1107 125 1109 129
rect 1113 125 1115 129
rect 1119 125 1121 129
rect 1125 125 1127 129
rect 1131 125 1133 129
rect 1137 125 1139 129
rect 1103 123 1143 125
rect 1107 119 1109 123
rect 1113 119 1115 123
rect 1119 119 1121 123
rect 1125 119 1127 123
rect 1131 119 1133 123
rect 1137 119 1139 123
rect 1103 116 1143 119
rect 1107 112 1109 116
rect 1113 112 1115 116
rect 1119 112 1121 116
rect 1125 112 1127 116
rect 1131 112 1133 116
rect 1137 112 1139 116
rect 1103 111 1143 112
rect 1107 107 1109 111
rect 1113 107 1115 111
rect 1119 107 1121 111
rect 1125 107 1127 111
rect 1131 107 1133 111
rect 1137 107 1139 111
rect 973 92 975 101
rect 979 92 981 101
rect 985 92 987 101
rect 991 92 993 101
rect 997 92 999 101
rect 1003 92 1005 101
rect 1147 101 1187 137
rect 969 90 1009 92
rect 973 86 975 90
rect 979 86 981 90
rect 985 86 987 90
rect 991 86 993 90
rect 997 86 999 90
rect 1003 86 1005 90
rect 969 84 1009 86
rect 973 80 975 84
rect 979 80 981 84
rect 985 80 987 84
rect 991 80 993 84
rect 997 80 999 84
rect 1003 80 1005 84
rect 969 78 1009 80
rect 973 74 975 78
rect 979 74 981 78
rect 985 74 987 78
rect 991 74 993 78
rect 997 74 999 78
rect 1003 74 1005 78
rect 969 72 1009 74
rect 973 63 975 72
rect 979 63 981 72
rect 985 63 987 72
rect 991 63 993 72
rect 997 63 999 72
rect 1003 63 1005 72
rect 969 12 1009 63
rect 973 8 975 12
rect 979 8 981 12
rect 985 8 987 12
rect 991 8 993 12
rect 997 8 999 12
rect 1003 8 1005 12
rect 969 4 1009 8
rect 973 0 975 4
rect 979 0 981 4
rect 985 0 987 4
rect 991 0 993 4
rect 997 0 999 4
rect 1003 0 1005 4
rect 1013 99 1043 100
rect 1013 95 1014 99
rect 1018 95 1020 99
rect 1024 95 1026 99
rect 1030 95 1032 99
rect 1036 95 1038 99
rect 1042 95 1043 99
rect 1013 93 1043 95
rect 1013 89 1014 93
rect 1018 89 1020 93
rect 1024 89 1026 93
rect 1030 89 1032 93
rect 1036 89 1038 93
rect 1042 89 1043 93
rect 1013 86 1043 89
rect 1013 82 1014 86
rect 1018 82 1020 86
rect 1024 82 1026 86
rect 1030 82 1032 86
rect 1036 82 1038 86
rect 1042 82 1043 86
rect 1013 80 1043 82
rect 1013 76 1014 80
rect 1018 76 1020 80
rect 1024 76 1026 80
rect 1030 76 1032 80
rect 1036 76 1038 80
rect 1042 76 1043 80
rect 1013 74 1043 76
rect 1013 70 1014 74
rect 1018 70 1020 74
rect 1024 70 1026 74
rect 1030 70 1032 74
rect 1036 70 1038 74
rect 1042 70 1043 74
rect 1013 68 1043 70
rect 1013 64 1014 68
rect 1018 64 1020 68
rect 1024 64 1026 68
rect 1030 64 1032 68
rect 1036 64 1038 68
rect 1042 64 1043 68
rect 1013 48 1043 64
rect 1113 99 1143 100
rect 1113 95 1114 99
rect 1118 95 1120 99
rect 1124 95 1126 99
rect 1130 95 1132 99
rect 1136 95 1138 99
rect 1142 95 1143 99
rect 1113 93 1143 95
rect 1113 89 1114 93
rect 1118 89 1120 93
rect 1124 89 1126 93
rect 1130 89 1132 93
rect 1136 89 1138 93
rect 1142 89 1143 93
rect 1113 86 1143 89
rect 1113 82 1114 86
rect 1118 82 1120 86
rect 1124 82 1126 86
rect 1130 82 1132 86
rect 1136 82 1138 86
rect 1142 82 1143 86
rect 1113 80 1143 82
rect 1113 76 1114 80
rect 1118 76 1120 80
rect 1124 76 1126 80
rect 1130 76 1132 80
rect 1136 76 1138 80
rect 1142 76 1143 80
rect 1113 74 1143 76
rect 1113 70 1114 74
rect 1118 70 1120 74
rect 1124 70 1126 74
rect 1130 70 1132 74
rect 1136 70 1138 74
rect 1142 70 1143 74
rect 1113 68 1143 70
rect 1113 64 1114 68
rect 1118 64 1120 68
rect 1124 64 1126 68
rect 1130 64 1132 68
rect 1136 64 1138 68
rect 1142 64 1143 68
rect 1047 57 1066 58
rect 1051 53 1052 57
rect 1056 53 1057 57
rect 1061 53 1062 57
rect 1047 52 1066 53
rect 1017 44 1019 48
rect 1023 44 1025 48
rect 1029 44 1031 48
rect 1035 44 1037 48
rect 1041 44 1043 48
rect 1047 44 1049 48
rect 1013 42 1053 44
rect 1017 38 1019 42
rect 1023 38 1025 42
rect 1029 38 1031 42
rect 1035 38 1037 42
rect 1041 38 1043 42
rect 1047 38 1049 42
rect 1013 36 1053 38
rect 1017 32 1019 36
rect 1023 32 1025 36
rect 1029 32 1031 36
rect 1035 32 1037 36
rect 1041 32 1043 36
rect 1047 32 1049 36
rect 1013 30 1053 32
rect 1017 26 1019 30
rect 1023 26 1025 30
rect 1029 26 1031 30
rect 1035 26 1037 30
rect 1041 26 1043 30
rect 1047 26 1049 30
rect 1013 24 1053 26
rect 1017 20 1019 24
rect 1023 20 1025 24
rect 1029 20 1031 24
rect 1035 20 1037 24
rect 1041 20 1043 24
rect 1047 20 1049 24
rect 1013 18 1053 20
rect 1013 14 1019 18
rect 1023 14 1025 18
rect 1029 14 1031 18
rect 1035 14 1037 18
rect 1041 14 1043 18
rect 1047 14 1049 18
rect 1013 4 1053 14
rect 1017 0 1019 4
rect 1023 0 1025 4
rect 1029 0 1031 4
rect 1035 0 1037 4
rect 1041 0 1043 4
rect 1047 0 1049 4
rect 1057 4 1066 52
rect 1090 57 1109 58
rect 1094 53 1095 57
rect 1099 53 1100 57
rect 1104 53 1105 57
rect 1090 52 1109 53
rect 1090 4 1099 52
rect 1113 48 1143 64
rect 1107 44 1109 48
rect 1113 44 1115 48
rect 1119 44 1121 48
rect 1125 44 1127 48
rect 1131 44 1133 48
rect 1137 44 1139 48
rect 1103 42 1143 44
rect 1107 38 1109 42
rect 1113 38 1115 42
rect 1119 38 1121 42
rect 1125 38 1127 42
rect 1131 38 1133 42
rect 1137 38 1139 42
rect 1103 36 1143 38
rect 1107 32 1109 36
rect 1113 32 1115 36
rect 1119 32 1121 36
rect 1125 32 1127 36
rect 1131 32 1133 36
rect 1137 32 1139 36
rect 1103 30 1143 32
rect 1107 26 1109 30
rect 1113 26 1115 30
rect 1119 26 1121 30
rect 1125 26 1127 30
rect 1131 26 1133 30
rect 1137 26 1139 30
rect 1103 24 1143 26
rect 1107 20 1109 24
rect 1113 20 1115 24
rect 1119 20 1121 24
rect 1125 20 1127 24
rect 1131 20 1133 24
rect 1137 20 1139 24
rect 1103 18 1143 20
rect 1107 14 1109 18
rect 1113 14 1115 18
rect 1119 14 1121 18
rect 1125 14 1127 18
rect 1131 14 1133 18
rect 1137 14 1143 18
rect 1103 4 1143 14
rect 1107 0 1109 4
rect 1113 0 1115 4
rect 1119 0 1121 4
rect 1125 0 1127 4
rect 1131 0 1133 4
rect 1137 0 1139 4
rect 1151 92 1153 101
rect 1157 92 1159 101
rect 1163 92 1165 101
rect 1169 92 1171 101
rect 1175 92 1177 101
rect 1181 92 1183 101
rect 1147 90 1187 92
rect 1151 86 1153 90
rect 1157 86 1159 90
rect 1163 86 1165 90
rect 1169 86 1171 90
rect 1175 86 1177 90
rect 1181 86 1183 90
rect 1147 84 1187 86
rect 1151 80 1153 84
rect 1157 80 1159 84
rect 1163 80 1165 84
rect 1169 80 1171 84
rect 1175 80 1177 84
rect 1181 80 1183 84
rect 1147 78 1187 80
rect 1151 74 1153 78
rect 1157 74 1159 78
rect 1163 74 1165 78
rect 1169 74 1171 78
rect 1175 74 1177 78
rect 1181 74 1183 78
rect 1147 72 1187 74
rect 1151 63 1153 72
rect 1157 63 1159 72
rect 1163 63 1165 72
rect 1169 63 1171 72
rect 1175 63 1177 72
rect 1181 63 1183 72
rect 1147 12 1187 63
rect 1151 8 1153 12
rect 1157 8 1159 12
rect 1163 8 1165 12
rect 1169 8 1171 12
rect 1175 8 1177 12
rect 1181 8 1183 12
rect 1147 4 1187 8
rect 1151 0 1153 4
rect 1157 0 1159 4
rect 1163 0 1165 4
rect 1169 0 1171 4
rect 1175 0 1177 4
rect 1181 0 1183 4
rect 1443 141 1483 144
rect 1447 137 1449 141
rect 1453 137 1455 141
rect 1459 137 1461 141
rect 1465 137 1467 141
rect 1471 137 1473 141
rect 1477 137 1479 141
rect 1443 101 1483 137
rect 1621 141 1661 144
rect 1625 137 1627 141
rect 1631 137 1633 141
rect 1637 137 1639 141
rect 1643 137 1645 141
rect 1649 137 1651 141
rect 1655 137 1657 141
rect 1497 131 1499 135
rect 1503 131 1505 135
rect 1509 131 1511 135
rect 1515 131 1517 135
rect 1521 131 1523 135
rect 1493 129 1527 131
rect 1491 125 1493 129
rect 1497 125 1499 129
rect 1503 125 1505 129
rect 1509 125 1511 129
rect 1515 125 1517 129
rect 1521 125 1523 129
rect 1487 123 1527 125
rect 1491 119 1493 123
rect 1497 119 1499 123
rect 1503 119 1505 123
rect 1509 119 1511 123
rect 1515 119 1517 123
rect 1521 119 1523 123
rect 1487 116 1527 119
rect 1491 112 1493 116
rect 1497 112 1499 116
rect 1503 112 1505 116
rect 1509 112 1511 116
rect 1515 112 1517 116
rect 1521 112 1523 116
rect 1487 111 1527 112
rect 1491 107 1493 111
rect 1497 107 1499 111
rect 1503 107 1505 111
rect 1509 107 1511 111
rect 1515 107 1517 111
rect 1521 107 1523 111
rect 1581 131 1583 135
rect 1587 131 1589 135
rect 1593 131 1595 135
rect 1599 131 1601 135
rect 1605 131 1607 135
rect 1577 129 1611 131
rect 1581 125 1583 129
rect 1587 125 1589 129
rect 1593 125 1595 129
rect 1599 125 1601 129
rect 1605 125 1607 129
rect 1611 125 1613 129
rect 1577 123 1617 125
rect 1581 119 1583 123
rect 1587 119 1589 123
rect 1593 119 1595 123
rect 1599 119 1601 123
rect 1605 119 1607 123
rect 1611 119 1613 123
rect 1577 116 1617 119
rect 1581 112 1583 116
rect 1587 112 1589 116
rect 1593 112 1595 116
rect 1599 112 1601 116
rect 1605 112 1607 116
rect 1611 112 1613 116
rect 1577 111 1617 112
rect 1581 107 1583 111
rect 1587 107 1589 111
rect 1593 107 1595 111
rect 1599 107 1601 111
rect 1605 107 1607 111
rect 1611 107 1613 111
rect 1447 92 1449 101
rect 1453 92 1455 101
rect 1459 92 1461 101
rect 1465 92 1467 101
rect 1471 92 1473 101
rect 1477 92 1479 101
rect 1621 101 1661 137
rect 1443 90 1483 92
rect 1447 86 1449 90
rect 1453 86 1455 90
rect 1459 86 1461 90
rect 1465 86 1467 90
rect 1471 86 1473 90
rect 1477 86 1479 90
rect 1443 84 1483 86
rect 1447 80 1449 84
rect 1453 80 1455 84
rect 1459 80 1461 84
rect 1465 80 1467 84
rect 1471 80 1473 84
rect 1477 80 1479 84
rect 1443 78 1483 80
rect 1447 74 1449 78
rect 1453 74 1455 78
rect 1459 74 1461 78
rect 1465 74 1467 78
rect 1471 74 1473 78
rect 1477 74 1479 78
rect 1443 72 1483 74
rect 1447 63 1449 72
rect 1453 63 1455 72
rect 1459 63 1461 72
rect 1465 63 1467 72
rect 1471 63 1473 72
rect 1477 63 1479 72
rect 1443 12 1483 63
rect 1447 8 1449 12
rect 1453 8 1455 12
rect 1459 8 1461 12
rect 1465 8 1467 12
rect 1471 8 1473 12
rect 1477 8 1479 12
rect 1443 4 1483 8
rect 1447 0 1449 4
rect 1453 0 1455 4
rect 1459 0 1461 4
rect 1465 0 1467 4
rect 1471 0 1473 4
rect 1477 0 1479 4
rect 1487 99 1517 100
rect 1487 95 1488 99
rect 1492 95 1494 99
rect 1498 95 1500 99
rect 1504 95 1506 99
rect 1510 95 1512 99
rect 1516 95 1517 99
rect 1487 93 1517 95
rect 1487 89 1488 93
rect 1492 89 1494 93
rect 1498 89 1500 93
rect 1504 89 1506 93
rect 1510 89 1512 93
rect 1516 89 1517 93
rect 1487 86 1517 89
rect 1487 82 1488 86
rect 1492 82 1494 86
rect 1498 82 1500 86
rect 1504 82 1506 86
rect 1510 82 1512 86
rect 1516 82 1517 86
rect 1487 80 1517 82
rect 1487 76 1488 80
rect 1492 76 1494 80
rect 1498 76 1500 80
rect 1504 76 1506 80
rect 1510 76 1512 80
rect 1516 76 1517 80
rect 1487 74 1517 76
rect 1487 70 1488 74
rect 1492 70 1494 74
rect 1498 70 1500 74
rect 1504 70 1506 74
rect 1510 70 1512 74
rect 1516 70 1517 74
rect 1487 68 1517 70
rect 1487 64 1488 68
rect 1492 64 1494 68
rect 1498 64 1500 68
rect 1504 64 1506 68
rect 1510 64 1512 68
rect 1516 64 1517 68
rect 1487 48 1517 64
rect 1587 99 1617 100
rect 1587 95 1588 99
rect 1592 95 1594 99
rect 1598 95 1600 99
rect 1604 95 1606 99
rect 1610 95 1612 99
rect 1616 95 1617 99
rect 1587 93 1617 95
rect 1587 89 1588 93
rect 1592 89 1594 93
rect 1598 89 1600 93
rect 1604 89 1606 93
rect 1610 89 1612 93
rect 1616 89 1617 93
rect 1587 86 1617 89
rect 1587 82 1588 86
rect 1592 82 1594 86
rect 1598 82 1600 86
rect 1604 82 1606 86
rect 1610 82 1612 86
rect 1616 82 1617 86
rect 1587 80 1617 82
rect 1587 76 1588 80
rect 1592 76 1594 80
rect 1598 76 1600 80
rect 1604 76 1606 80
rect 1610 76 1612 80
rect 1616 76 1617 80
rect 1587 74 1617 76
rect 1587 70 1588 74
rect 1592 70 1594 74
rect 1598 70 1600 74
rect 1604 70 1606 74
rect 1610 70 1612 74
rect 1616 70 1617 74
rect 1587 68 1617 70
rect 1587 64 1588 68
rect 1592 64 1594 68
rect 1598 64 1600 68
rect 1604 64 1606 68
rect 1610 64 1612 68
rect 1616 64 1617 68
rect 1521 57 1540 58
rect 1525 53 1526 57
rect 1530 53 1531 57
rect 1535 53 1536 57
rect 1521 52 1540 53
rect 1491 44 1493 48
rect 1497 44 1499 48
rect 1503 44 1505 48
rect 1509 44 1511 48
rect 1515 44 1517 48
rect 1521 44 1523 48
rect 1487 42 1527 44
rect 1491 38 1493 42
rect 1497 38 1499 42
rect 1503 38 1505 42
rect 1509 38 1511 42
rect 1515 38 1517 42
rect 1521 38 1523 42
rect 1487 36 1527 38
rect 1491 32 1493 36
rect 1497 32 1499 36
rect 1503 32 1505 36
rect 1509 32 1511 36
rect 1515 32 1517 36
rect 1521 32 1523 36
rect 1487 30 1527 32
rect 1491 26 1493 30
rect 1497 26 1499 30
rect 1503 26 1505 30
rect 1509 26 1511 30
rect 1515 26 1517 30
rect 1521 26 1523 30
rect 1487 24 1527 26
rect 1491 20 1493 24
rect 1497 20 1499 24
rect 1503 20 1505 24
rect 1509 20 1511 24
rect 1515 20 1517 24
rect 1521 20 1523 24
rect 1487 18 1527 20
rect 1487 14 1493 18
rect 1497 14 1499 18
rect 1503 14 1505 18
rect 1509 14 1511 18
rect 1515 14 1517 18
rect 1521 14 1523 18
rect 1487 4 1527 14
rect 1491 0 1493 4
rect 1497 0 1499 4
rect 1503 0 1505 4
rect 1509 0 1511 4
rect 1515 0 1517 4
rect 1521 0 1523 4
rect 1531 4 1540 52
rect 1564 57 1583 58
rect 1568 53 1569 57
rect 1573 53 1574 57
rect 1578 53 1579 57
rect 1564 52 1583 53
rect 1564 4 1573 52
rect 1587 48 1617 64
rect 1581 44 1583 48
rect 1587 44 1589 48
rect 1593 44 1595 48
rect 1599 44 1601 48
rect 1605 44 1607 48
rect 1611 44 1613 48
rect 1577 42 1617 44
rect 1581 38 1583 42
rect 1587 38 1589 42
rect 1593 38 1595 42
rect 1599 38 1601 42
rect 1605 38 1607 42
rect 1611 38 1613 42
rect 1577 36 1617 38
rect 1581 32 1583 36
rect 1587 32 1589 36
rect 1593 32 1595 36
rect 1599 32 1601 36
rect 1605 32 1607 36
rect 1611 32 1613 36
rect 1577 30 1617 32
rect 1581 26 1583 30
rect 1587 26 1589 30
rect 1593 26 1595 30
rect 1599 26 1601 30
rect 1605 26 1607 30
rect 1611 26 1613 30
rect 1577 24 1617 26
rect 1581 20 1583 24
rect 1587 20 1589 24
rect 1593 20 1595 24
rect 1599 20 1601 24
rect 1605 20 1607 24
rect 1611 20 1613 24
rect 1577 18 1617 20
rect 1581 14 1583 18
rect 1587 14 1589 18
rect 1593 14 1595 18
rect 1599 14 1601 18
rect 1605 14 1607 18
rect 1611 14 1617 18
rect 1577 4 1617 14
rect 1581 0 1583 4
rect 1587 0 1589 4
rect 1593 0 1595 4
rect 1599 0 1601 4
rect 1605 0 1607 4
rect 1611 0 1613 4
rect 1625 92 1627 101
rect 1631 92 1633 101
rect 1637 92 1639 101
rect 1643 92 1645 101
rect 1649 92 1651 101
rect 1655 92 1657 101
rect 1621 90 1661 92
rect 1625 86 1627 90
rect 1631 86 1633 90
rect 1637 86 1639 90
rect 1643 86 1645 90
rect 1649 86 1651 90
rect 1655 86 1657 90
rect 1621 84 1661 86
rect 1625 80 1627 84
rect 1631 80 1633 84
rect 1637 80 1639 84
rect 1643 80 1645 84
rect 1649 80 1651 84
rect 1655 80 1657 84
rect 1621 78 1661 80
rect 1625 74 1627 78
rect 1631 74 1633 78
rect 1637 74 1639 78
rect 1643 74 1645 78
rect 1649 74 1651 78
rect 1655 74 1657 78
rect 1621 72 1661 74
rect 1625 63 1627 72
rect 1631 63 1633 72
rect 1637 63 1639 72
rect 1643 63 1645 72
rect 1649 63 1651 72
rect 1655 63 1657 72
rect 1621 12 1661 63
rect 1625 8 1627 12
rect 1631 8 1633 12
rect 1637 8 1639 12
rect 1643 8 1645 12
rect 1649 8 1651 12
rect 1655 8 1657 12
rect 1621 4 1661 8
rect 1625 0 1627 4
rect 1631 0 1633 4
rect 1637 0 1639 4
rect 1643 0 1645 4
rect 1649 0 1651 4
rect 1655 0 1657 4
rect 1917 141 1957 144
rect 1921 137 1923 141
rect 1927 137 1929 141
rect 1933 137 1935 141
rect 1939 137 1941 141
rect 1945 137 1947 141
rect 1951 137 1953 141
rect 1917 101 1957 137
rect 2095 141 2135 144
rect 2099 137 2101 141
rect 2105 137 2107 141
rect 2111 137 2113 141
rect 2117 137 2119 141
rect 2123 137 2125 141
rect 2129 137 2131 141
rect 1971 131 1973 135
rect 1977 131 1979 135
rect 1983 131 1985 135
rect 1989 131 1991 135
rect 1995 131 1997 135
rect 1967 129 2001 131
rect 1965 125 1967 129
rect 1971 125 1973 129
rect 1977 125 1979 129
rect 1983 125 1985 129
rect 1989 125 1991 129
rect 1995 125 1997 129
rect 1961 123 2001 125
rect 1965 119 1967 123
rect 1971 119 1973 123
rect 1977 119 1979 123
rect 1983 119 1985 123
rect 1989 119 1991 123
rect 1995 119 1997 123
rect 1961 116 2001 119
rect 1965 112 1967 116
rect 1971 112 1973 116
rect 1977 112 1979 116
rect 1983 112 1985 116
rect 1989 112 1991 116
rect 1995 112 1997 116
rect 1961 111 2001 112
rect 1965 107 1967 111
rect 1971 107 1973 111
rect 1977 107 1979 111
rect 1983 107 1985 111
rect 1989 107 1991 111
rect 1995 107 1997 111
rect 2055 131 2057 135
rect 2061 131 2063 135
rect 2067 131 2069 135
rect 2073 131 2075 135
rect 2079 131 2081 135
rect 2051 129 2085 131
rect 2055 125 2057 129
rect 2061 125 2063 129
rect 2067 125 2069 129
rect 2073 125 2075 129
rect 2079 125 2081 129
rect 2085 125 2087 129
rect 2051 123 2091 125
rect 2055 119 2057 123
rect 2061 119 2063 123
rect 2067 119 2069 123
rect 2073 119 2075 123
rect 2079 119 2081 123
rect 2085 119 2087 123
rect 2051 116 2091 119
rect 2055 112 2057 116
rect 2061 112 2063 116
rect 2067 112 2069 116
rect 2073 112 2075 116
rect 2079 112 2081 116
rect 2085 112 2087 116
rect 2051 111 2091 112
rect 2055 107 2057 111
rect 2061 107 2063 111
rect 2067 107 2069 111
rect 2073 107 2075 111
rect 2079 107 2081 111
rect 2085 107 2087 111
rect 1921 92 1923 101
rect 1927 92 1929 101
rect 1933 92 1935 101
rect 1939 92 1941 101
rect 1945 92 1947 101
rect 1951 92 1953 101
rect 2095 101 2135 137
rect 1917 90 1957 92
rect 1921 86 1923 90
rect 1927 86 1929 90
rect 1933 86 1935 90
rect 1939 86 1941 90
rect 1945 86 1947 90
rect 1951 86 1953 90
rect 1917 84 1957 86
rect 1921 80 1923 84
rect 1927 80 1929 84
rect 1933 80 1935 84
rect 1939 80 1941 84
rect 1945 80 1947 84
rect 1951 80 1953 84
rect 1917 78 1957 80
rect 1921 74 1923 78
rect 1927 74 1929 78
rect 1933 74 1935 78
rect 1939 74 1941 78
rect 1945 74 1947 78
rect 1951 74 1953 78
rect 1917 72 1957 74
rect 1921 63 1923 72
rect 1927 63 1929 72
rect 1933 63 1935 72
rect 1939 63 1941 72
rect 1945 63 1947 72
rect 1951 63 1953 72
rect 1917 12 1957 63
rect 1921 8 1923 12
rect 1927 8 1929 12
rect 1933 8 1935 12
rect 1939 8 1941 12
rect 1945 8 1947 12
rect 1951 8 1953 12
rect 1917 4 1957 8
rect 1921 0 1923 4
rect 1927 0 1929 4
rect 1933 0 1935 4
rect 1939 0 1941 4
rect 1945 0 1947 4
rect 1951 0 1953 4
rect 1961 99 1991 100
rect 1961 95 1962 99
rect 1966 95 1968 99
rect 1972 95 1974 99
rect 1978 95 1980 99
rect 1984 95 1986 99
rect 1990 95 1991 99
rect 1961 93 1991 95
rect 1961 89 1962 93
rect 1966 89 1968 93
rect 1972 89 1974 93
rect 1978 89 1980 93
rect 1984 89 1986 93
rect 1990 89 1991 93
rect 1961 86 1991 89
rect 1961 82 1962 86
rect 1966 82 1968 86
rect 1972 82 1974 86
rect 1978 82 1980 86
rect 1984 82 1986 86
rect 1990 82 1991 86
rect 1961 80 1991 82
rect 1961 76 1962 80
rect 1966 76 1968 80
rect 1972 76 1974 80
rect 1978 76 1980 80
rect 1984 76 1986 80
rect 1990 76 1991 80
rect 1961 74 1991 76
rect 1961 70 1962 74
rect 1966 70 1968 74
rect 1972 70 1974 74
rect 1978 70 1980 74
rect 1984 70 1986 74
rect 1990 70 1991 74
rect 1961 68 1991 70
rect 1961 64 1962 68
rect 1966 64 1968 68
rect 1972 64 1974 68
rect 1978 64 1980 68
rect 1984 64 1986 68
rect 1990 64 1991 68
rect 1961 48 1991 64
rect 2061 99 2091 100
rect 2061 95 2062 99
rect 2066 95 2068 99
rect 2072 95 2074 99
rect 2078 95 2080 99
rect 2084 95 2086 99
rect 2090 95 2091 99
rect 2061 93 2091 95
rect 2061 89 2062 93
rect 2066 89 2068 93
rect 2072 89 2074 93
rect 2078 89 2080 93
rect 2084 89 2086 93
rect 2090 89 2091 93
rect 2061 86 2091 89
rect 2061 82 2062 86
rect 2066 82 2068 86
rect 2072 82 2074 86
rect 2078 82 2080 86
rect 2084 82 2086 86
rect 2090 82 2091 86
rect 2061 80 2091 82
rect 2061 76 2062 80
rect 2066 76 2068 80
rect 2072 76 2074 80
rect 2078 76 2080 80
rect 2084 76 2086 80
rect 2090 76 2091 80
rect 2061 74 2091 76
rect 2061 70 2062 74
rect 2066 70 2068 74
rect 2072 70 2074 74
rect 2078 70 2080 74
rect 2084 70 2086 74
rect 2090 70 2091 74
rect 2061 68 2091 70
rect 2061 64 2062 68
rect 2066 64 2068 68
rect 2072 64 2074 68
rect 2078 64 2080 68
rect 2084 64 2086 68
rect 2090 64 2091 68
rect 1995 57 2014 58
rect 1999 53 2000 57
rect 2004 53 2005 57
rect 2009 53 2010 57
rect 1995 52 2014 53
rect 1965 44 1967 48
rect 1971 44 1973 48
rect 1977 44 1979 48
rect 1983 44 1985 48
rect 1989 44 1991 48
rect 1995 44 1997 48
rect 1961 42 2001 44
rect 1965 38 1967 42
rect 1971 38 1973 42
rect 1977 38 1979 42
rect 1983 38 1985 42
rect 1989 38 1991 42
rect 1995 38 1997 42
rect 1961 36 2001 38
rect 1965 32 1967 36
rect 1971 32 1973 36
rect 1977 32 1979 36
rect 1983 32 1985 36
rect 1989 32 1991 36
rect 1995 32 1997 36
rect 1961 30 2001 32
rect 1965 26 1967 30
rect 1971 26 1973 30
rect 1977 26 1979 30
rect 1983 26 1985 30
rect 1989 26 1991 30
rect 1995 26 1997 30
rect 1961 24 2001 26
rect 1965 20 1967 24
rect 1971 20 1973 24
rect 1977 20 1979 24
rect 1983 20 1985 24
rect 1989 20 1991 24
rect 1995 20 1997 24
rect 1961 18 2001 20
rect 1961 14 1967 18
rect 1971 14 1973 18
rect 1977 14 1979 18
rect 1983 14 1985 18
rect 1989 14 1991 18
rect 1995 14 1997 18
rect 1961 4 2001 14
rect 1965 0 1967 4
rect 1971 0 1973 4
rect 1977 0 1979 4
rect 1983 0 1985 4
rect 1989 0 1991 4
rect 1995 0 1997 4
rect 2005 4 2014 52
rect 2038 57 2057 58
rect 2042 53 2043 57
rect 2047 53 2048 57
rect 2052 53 2053 57
rect 2038 52 2057 53
rect 2038 4 2047 52
rect 2061 48 2091 64
rect 2055 44 2057 48
rect 2061 44 2063 48
rect 2067 44 2069 48
rect 2073 44 2075 48
rect 2079 44 2081 48
rect 2085 44 2087 48
rect 2051 42 2091 44
rect 2055 38 2057 42
rect 2061 38 2063 42
rect 2067 38 2069 42
rect 2073 38 2075 42
rect 2079 38 2081 42
rect 2085 38 2087 42
rect 2051 36 2091 38
rect 2055 32 2057 36
rect 2061 32 2063 36
rect 2067 32 2069 36
rect 2073 32 2075 36
rect 2079 32 2081 36
rect 2085 32 2087 36
rect 2051 30 2091 32
rect 2055 26 2057 30
rect 2061 26 2063 30
rect 2067 26 2069 30
rect 2073 26 2075 30
rect 2079 26 2081 30
rect 2085 26 2087 30
rect 2051 24 2091 26
rect 2055 20 2057 24
rect 2061 20 2063 24
rect 2067 20 2069 24
rect 2073 20 2075 24
rect 2079 20 2081 24
rect 2085 20 2087 24
rect 2051 18 2091 20
rect 2055 14 2057 18
rect 2061 14 2063 18
rect 2067 14 2069 18
rect 2073 14 2075 18
rect 2079 14 2081 18
rect 2085 14 2091 18
rect 2051 4 2091 14
rect 2055 0 2057 4
rect 2061 0 2063 4
rect 2067 0 2069 4
rect 2073 0 2075 4
rect 2079 0 2081 4
rect 2085 0 2087 4
rect 2099 92 2101 101
rect 2105 92 2107 101
rect 2111 92 2113 101
rect 2117 92 2119 101
rect 2123 92 2125 101
rect 2129 92 2131 101
rect 2095 90 2135 92
rect 2099 86 2101 90
rect 2105 86 2107 90
rect 2111 86 2113 90
rect 2117 86 2119 90
rect 2123 86 2125 90
rect 2129 86 2131 90
rect 2095 84 2135 86
rect 2099 80 2101 84
rect 2105 80 2107 84
rect 2111 80 2113 84
rect 2117 80 2119 84
rect 2123 80 2125 84
rect 2129 80 2131 84
rect 2095 78 2135 80
rect 2099 74 2101 78
rect 2105 74 2107 78
rect 2111 74 2113 78
rect 2117 74 2119 78
rect 2123 74 2125 78
rect 2129 74 2131 78
rect 2095 72 2135 74
rect 2099 63 2101 72
rect 2105 63 2107 72
rect 2111 63 2113 72
rect 2117 63 2119 72
rect 2123 63 2125 72
rect 2129 63 2131 72
rect 2095 12 2135 63
rect 2099 8 2101 12
rect 2105 8 2107 12
rect 2111 8 2113 12
rect 2117 8 2119 12
rect 2123 8 2125 12
rect 2129 8 2131 12
rect 2095 4 2135 8
rect 2099 0 2101 4
rect 2105 0 2107 4
rect 2111 0 2113 4
rect 2117 0 2119 4
rect 2123 0 2125 4
rect 2129 0 2131 4
rect 2391 141 2431 144
rect 2395 137 2397 141
rect 2401 137 2403 141
rect 2407 137 2409 141
rect 2413 137 2415 141
rect 2419 137 2421 141
rect 2425 137 2427 141
rect 2391 101 2431 137
rect 2569 141 2609 144
rect 2573 137 2575 141
rect 2579 137 2581 141
rect 2585 137 2587 141
rect 2591 137 2593 141
rect 2597 137 2599 141
rect 2603 137 2605 141
rect 2445 131 2447 135
rect 2451 131 2453 135
rect 2457 131 2459 135
rect 2463 131 2465 135
rect 2469 131 2471 135
rect 2441 129 2475 131
rect 2439 125 2441 129
rect 2445 125 2447 129
rect 2451 125 2453 129
rect 2457 125 2459 129
rect 2463 125 2465 129
rect 2469 125 2471 129
rect 2435 123 2475 125
rect 2439 119 2441 123
rect 2445 119 2447 123
rect 2451 119 2453 123
rect 2457 119 2459 123
rect 2463 119 2465 123
rect 2469 119 2471 123
rect 2435 116 2475 119
rect 2439 112 2441 116
rect 2445 112 2447 116
rect 2451 112 2453 116
rect 2457 112 2459 116
rect 2463 112 2465 116
rect 2469 112 2471 116
rect 2435 111 2475 112
rect 2439 107 2441 111
rect 2445 107 2447 111
rect 2451 107 2453 111
rect 2457 107 2459 111
rect 2463 107 2465 111
rect 2469 107 2471 111
rect 2529 131 2531 135
rect 2535 131 2537 135
rect 2541 131 2543 135
rect 2547 131 2549 135
rect 2553 131 2555 135
rect 2525 129 2559 131
rect 2529 125 2531 129
rect 2535 125 2537 129
rect 2541 125 2543 129
rect 2547 125 2549 129
rect 2553 125 2555 129
rect 2559 125 2561 129
rect 2525 123 2565 125
rect 2529 119 2531 123
rect 2535 119 2537 123
rect 2541 119 2543 123
rect 2547 119 2549 123
rect 2553 119 2555 123
rect 2559 119 2561 123
rect 2525 116 2565 119
rect 2529 112 2531 116
rect 2535 112 2537 116
rect 2541 112 2543 116
rect 2547 112 2549 116
rect 2553 112 2555 116
rect 2559 112 2561 116
rect 2525 111 2565 112
rect 2529 107 2531 111
rect 2535 107 2537 111
rect 2541 107 2543 111
rect 2547 107 2549 111
rect 2553 107 2555 111
rect 2559 107 2561 111
rect 2395 92 2397 101
rect 2401 92 2403 101
rect 2407 92 2409 101
rect 2413 92 2415 101
rect 2419 92 2421 101
rect 2425 92 2427 101
rect 2569 101 2609 137
rect 2391 90 2431 92
rect 2395 86 2397 90
rect 2401 86 2403 90
rect 2407 86 2409 90
rect 2413 86 2415 90
rect 2419 86 2421 90
rect 2425 86 2427 90
rect 2391 84 2431 86
rect 2395 80 2397 84
rect 2401 80 2403 84
rect 2407 80 2409 84
rect 2413 80 2415 84
rect 2419 80 2421 84
rect 2425 80 2427 84
rect 2391 78 2431 80
rect 2395 74 2397 78
rect 2401 74 2403 78
rect 2407 74 2409 78
rect 2413 74 2415 78
rect 2419 74 2421 78
rect 2425 74 2427 78
rect 2391 72 2431 74
rect 2395 63 2397 72
rect 2401 63 2403 72
rect 2407 63 2409 72
rect 2413 63 2415 72
rect 2419 63 2421 72
rect 2425 63 2427 72
rect 2391 12 2431 63
rect 2395 8 2397 12
rect 2401 8 2403 12
rect 2407 8 2409 12
rect 2413 8 2415 12
rect 2419 8 2421 12
rect 2425 8 2427 12
rect 2391 4 2431 8
rect 2395 0 2397 4
rect 2401 0 2403 4
rect 2407 0 2409 4
rect 2413 0 2415 4
rect 2419 0 2421 4
rect 2425 0 2427 4
rect 2435 99 2465 100
rect 2435 95 2436 99
rect 2440 95 2442 99
rect 2446 95 2448 99
rect 2452 95 2454 99
rect 2458 95 2460 99
rect 2464 95 2465 99
rect 2435 93 2465 95
rect 2435 89 2436 93
rect 2440 89 2442 93
rect 2446 89 2448 93
rect 2452 89 2454 93
rect 2458 89 2460 93
rect 2464 89 2465 93
rect 2435 86 2465 89
rect 2435 82 2436 86
rect 2440 82 2442 86
rect 2446 82 2448 86
rect 2452 82 2454 86
rect 2458 82 2460 86
rect 2464 82 2465 86
rect 2435 80 2465 82
rect 2435 76 2436 80
rect 2440 76 2442 80
rect 2446 76 2448 80
rect 2452 76 2454 80
rect 2458 76 2460 80
rect 2464 76 2465 80
rect 2435 74 2465 76
rect 2435 70 2436 74
rect 2440 70 2442 74
rect 2446 70 2448 74
rect 2452 70 2454 74
rect 2458 70 2460 74
rect 2464 70 2465 74
rect 2435 68 2465 70
rect 2435 64 2436 68
rect 2440 64 2442 68
rect 2446 64 2448 68
rect 2452 64 2454 68
rect 2458 64 2460 68
rect 2464 64 2465 68
rect 2435 48 2465 64
rect 2535 99 2565 100
rect 2535 95 2536 99
rect 2540 95 2542 99
rect 2546 95 2548 99
rect 2552 95 2554 99
rect 2558 95 2560 99
rect 2564 95 2565 99
rect 2535 93 2565 95
rect 2535 89 2536 93
rect 2540 89 2542 93
rect 2546 89 2548 93
rect 2552 89 2554 93
rect 2558 89 2560 93
rect 2564 89 2565 93
rect 2535 86 2565 89
rect 2535 82 2536 86
rect 2540 82 2542 86
rect 2546 82 2548 86
rect 2552 82 2554 86
rect 2558 82 2560 86
rect 2564 82 2565 86
rect 2535 80 2565 82
rect 2535 76 2536 80
rect 2540 76 2542 80
rect 2546 76 2548 80
rect 2552 76 2554 80
rect 2558 76 2560 80
rect 2564 76 2565 80
rect 2535 74 2565 76
rect 2535 70 2536 74
rect 2540 70 2542 74
rect 2546 70 2548 74
rect 2552 70 2554 74
rect 2558 70 2560 74
rect 2564 70 2565 74
rect 2535 68 2565 70
rect 2535 64 2536 68
rect 2540 64 2542 68
rect 2546 64 2548 68
rect 2552 64 2554 68
rect 2558 64 2560 68
rect 2564 64 2565 68
rect 2469 57 2488 58
rect 2473 53 2474 57
rect 2478 53 2479 57
rect 2483 53 2484 57
rect 2469 52 2488 53
rect 2439 44 2441 48
rect 2445 44 2447 48
rect 2451 44 2453 48
rect 2457 44 2459 48
rect 2463 44 2465 48
rect 2469 44 2471 48
rect 2435 42 2475 44
rect 2439 38 2441 42
rect 2445 38 2447 42
rect 2451 38 2453 42
rect 2457 38 2459 42
rect 2463 38 2465 42
rect 2469 38 2471 42
rect 2435 36 2475 38
rect 2439 32 2441 36
rect 2445 32 2447 36
rect 2451 32 2453 36
rect 2457 32 2459 36
rect 2463 32 2465 36
rect 2469 32 2471 36
rect 2435 30 2475 32
rect 2439 26 2441 30
rect 2445 26 2447 30
rect 2451 26 2453 30
rect 2457 26 2459 30
rect 2463 26 2465 30
rect 2469 26 2471 30
rect 2435 24 2475 26
rect 2439 20 2441 24
rect 2445 20 2447 24
rect 2451 20 2453 24
rect 2457 20 2459 24
rect 2463 20 2465 24
rect 2469 20 2471 24
rect 2435 18 2475 20
rect 2435 14 2441 18
rect 2445 14 2447 18
rect 2451 14 2453 18
rect 2457 14 2459 18
rect 2463 14 2465 18
rect 2469 14 2471 18
rect 2435 4 2475 14
rect 2439 0 2441 4
rect 2445 0 2447 4
rect 2451 0 2453 4
rect 2457 0 2459 4
rect 2463 0 2465 4
rect 2469 0 2471 4
rect 2479 4 2488 52
rect 2512 57 2531 58
rect 2516 53 2517 57
rect 2521 53 2522 57
rect 2526 53 2527 57
rect 2512 52 2531 53
rect 2512 4 2521 52
rect 2535 48 2565 64
rect 2529 44 2531 48
rect 2535 44 2537 48
rect 2541 44 2543 48
rect 2547 44 2549 48
rect 2553 44 2555 48
rect 2559 44 2561 48
rect 2525 42 2565 44
rect 2529 38 2531 42
rect 2535 38 2537 42
rect 2541 38 2543 42
rect 2547 38 2549 42
rect 2553 38 2555 42
rect 2559 38 2561 42
rect 2525 36 2565 38
rect 2529 32 2531 36
rect 2535 32 2537 36
rect 2541 32 2543 36
rect 2547 32 2549 36
rect 2553 32 2555 36
rect 2559 32 2561 36
rect 2525 30 2565 32
rect 2529 26 2531 30
rect 2535 26 2537 30
rect 2541 26 2543 30
rect 2547 26 2549 30
rect 2553 26 2555 30
rect 2559 26 2561 30
rect 2525 24 2565 26
rect 2529 20 2531 24
rect 2535 20 2537 24
rect 2541 20 2543 24
rect 2547 20 2549 24
rect 2553 20 2555 24
rect 2559 20 2561 24
rect 2525 18 2565 20
rect 2529 14 2531 18
rect 2535 14 2537 18
rect 2541 14 2543 18
rect 2547 14 2549 18
rect 2553 14 2555 18
rect 2559 14 2565 18
rect 2525 4 2565 14
rect 2529 0 2531 4
rect 2535 0 2537 4
rect 2541 0 2543 4
rect 2547 0 2549 4
rect 2553 0 2555 4
rect 2559 0 2561 4
rect 2573 92 2575 101
rect 2579 92 2581 101
rect 2585 92 2587 101
rect 2591 92 2593 101
rect 2597 92 2599 101
rect 2603 92 2605 101
rect 2569 90 2609 92
rect 2573 86 2575 90
rect 2579 86 2581 90
rect 2585 86 2587 90
rect 2591 86 2593 90
rect 2597 86 2599 90
rect 2603 86 2605 90
rect 2569 84 2609 86
rect 2573 80 2575 84
rect 2579 80 2581 84
rect 2585 80 2587 84
rect 2591 80 2593 84
rect 2597 80 2599 84
rect 2603 80 2605 84
rect 2569 78 2609 80
rect 2573 74 2575 78
rect 2579 74 2581 78
rect 2585 74 2587 78
rect 2591 74 2593 78
rect 2597 74 2599 78
rect 2603 74 2605 78
rect 2569 72 2609 74
rect 2573 63 2575 72
rect 2579 63 2581 72
rect 2585 63 2587 72
rect 2591 63 2593 72
rect 2597 63 2599 72
rect 2603 63 2605 72
rect 2569 12 2609 63
rect 2573 8 2575 12
rect 2579 8 2581 12
rect 2585 8 2587 12
rect 2591 8 2593 12
rect 2597 8 2599 12
rect 2603 8 2605 12
rect 2569 4 2609 8
rect 2573 0 2575 4
rect 2579 0 2581 4
rect 2585 0 2587 4
rect 2591 0 2593 4
rect 2597 0 2599 4
rect 2603 0 2605 4
rect 2865 141 2905 144
rect 2869 137 2871 141
rect 2875 137 2877 141
rect 2881 137 2883 141
rect 2887 137 2889 141
rect 2893 137 2895 141
rect 2899 137 2901 141
rect 2865 101 2905 137
rect 3043 141 3083 144
rect 3047 137 3049 141
rect 3053 137 3055 141
rect 3059 137 3061 141
rect 3065 137 3067 141
rect 3071 137 3073 141
rect 3077 137 3079 141
rect 2919 131 2921 135
rect 2925 131 2927 135
rect 2931 131 2933 135
rect 2937 131 2939 135
rect 2943 131 2945 135
rect 2915 129 2949 131
rect 2913 125 2915 129
rect 2919 125 2921 129
rect 2925 125 2927 129
rect 2931 125 2933 129
rect 2937 125 2939 129
rect 2943 125 2945 129
rect 2909 123 2949 125
rect 2913 119 2915 123
rect 2919 119 2921 123
rect 2925 119 2927 123
rect 2931 119 2933 123
rect 2937 119 2939 123
rect 2943 119 2945 123
rect 2909 116 2949 119
rect 2913 112 2915 116
rect 2919 112 2921 116
rect 2925 112 2927 116
rect 2931 112 2933 116
rect 2937 112 2939 116
rect 2943 112 2945 116
rect 2909 111 2949 112
rect 2913 107 2915 111
rect 2919 107 2921 111
rect 2925 107 2927 111
rect 2931 107 2933 111
rect 2937 107 2939 111
rect 2943 107 2945 111
rect 3003 131 3005 135
rect 3009 131 3011 135
rect 3015 131 3017 135
rect 3021 131 3023 135
rect 3027 131 3029 135
rect 2999 129 3033 131
rect 3003 125 3005 129
rect 3009 125 3011 129
rect 3015 125 3017 129
rect 3021 125 3023 129
rect 3027 125 3029 129
rect 3033 125 3035 129
rect 2999 123 3039 125
rect 3003 119 3005 123
rect 3009 119 3011 123
rect 3015 119 3017 123
rect 3021 119 3023 123
rect 3027 119 3029 123
rect 3033 119 3035 123
rect 2999 116 3039 119
rect 3003 112 3005 116
rect 3009 112 3011 116
rect 3015 112 3017 116
rect 3021 112 3023 116
rect 3027 112 3029 116
rect 3033 112 3035 116
rect 2999 111 3039 112
rect 3003 107 3005 111
rect 3009 107 3011 111
rect 3015 107 3017 111
rect 3021 107 3023 111
rect 3027 107 3029 111
rect 3033 107 3035 111
rect 2869 92 2871 101
rect 2875 92 2877 101
rect 2881 92 2883 101
rect 2887 92 2889 101
rect 2893 92 2895 101
rect 2899 92 2901 101
rect 3043 101 3083 137
rect 2865 90 2905 92
rect 2869 86 2871 90
rect 2875 86 2877 90
rect 2881 86 2883 90
rect 2887 86 2889 90
rect 2893 86 2895 90
rect 2899 86 2901 90
rect 2865 84 2905 86
rect 2869 80 2871 84
rect 2875 80 2877 84
rect 2881 80 2883 84
rect 2887 80 2889 84
rect 2893 80 2895 84
rect 2899 80 2901 84
rect 2865 78 2905 80
rect 2869 74 2871 78
rect 2875 74 2877 78
rect 2881 74 2883 78
rect 2887 74 2889 78
rect 2893 74 2895 78
rect 2899 74 2901 78
rect 2865 72 2905 74
rect 2869 63 2871 72
rect 2875 63 2877 72
rect 2881 63 2883 72
rect 2887 63 2889 72
rect 2893 63 2895 72
rect 2899 63 2901 72
rect 2865 12 2905 63
rect 2869 8 2871 12
rect 2875 8 2877 12
rect 2881 8 2883 12
rect 2887 8 2889 12
rect 2893 8 2895 12
rect 2899 8 2901 12
rect 2865 4 2905 8
rect 2869 0 2871 4
rect 2875 0 2877 4
rect 2881 0 2883 4
rect 2887 0 2889 4
rect 2893 0 2895 4
rect 2899 0 2901 4
rect 2909 99 2939 100
rect 2909 95 2910 99
rect 2914 95 2916 99
rect 2920 95 2922 99
rect 2926 95 2928 99
rect 2932 95 2934 99
rect 2938 95 2939 99
rect 2909 93 2939 95
rect 2909 89 2910 93
rect 2914 89 2916 93
rect 2920 89 2922 93
rect 2926 89 2928 93
rect 2932 89 2934 93
rect 2938 89 2939 93
rect 2909 86 2939 89
rect 2909 82 2910 86
rect 2914 82 2916 86
rect 2920 82 2922 86
rect 2926 82 2928 86
rect 2932 82 2934 86
rect 2938 82 2939 86
rect 2909 80 2939 82
rect 2909 76 2910 80
rect 2914 76 2916 80
rect 2920 76 2922 80
rect 2926 76 2928 80
rect 2932 76 2934 80
rect 2938 76 2939 80
rect 2909 74 2939 76
rect 2909 70 2910 74
rect 2914 70 2916 74
rect 2920 70 2922 74
rect 2926 70 2928 74
rect 2932 70 2934 74
rect 2938 70 2939 74
rect 2909 68 2939 70
rect 2909 64 2910 68
rect 2914 64 2916 68
rect 2920 64 2922 68
rect 2926 64 2928 68
rect 2932 64 2934 68
rect 2938 64 2939 68
rect 2909 48 2939 64
rect 3009 99 3039 100
rect 3009 95 3010 99
rect 3014 95 3016 99
rect 3020 95 3022 99
rect 3026 95 3028 99
rect 3032 95 3034 99
rect 3038 95 3039 99
rect 3009 93 3039 95
rect 3009 89 3010 93
rect 3014 89 3016 93
rect 3020 89 3022 93
rect 3026 89 3028 93
rect 3032 89 3034 93
rect 3038 89 3039 93
rect 3009 86 3039 89
rect 3009 82 3010 86
rect 3014 82 3016 86
rect 3020 82 3022 86
rect 3026 82 3028 86
rect 3032 82 3034 86
rect 3038 82 3039 86
rect 3009 80 3039 82
rect 3009 76 3010 80
rect 3014 76 3016 80
rect 3020 76 3022 80
rect 3026 76 3028 80
rect 3032 76 3034 80
rect 3038 76 3039 80
rect 3009 74 3039 76
rect 3009 70 3010 74
rect 3014 70 3016 74
rect 3020 70 3022 74
rect 3026 70 3028 74
rect 3032 70 3034 74
rect 3038 70 3039 74
rect 3009 68 3039 70
rect 3009 64 3010 68
rect 3014 64 3016 68
rect 3020 64 3022 68
rect 3026 64 3028 68
rect 3032 64 3034 68
rect 3038 64 3039 68
rect 2943 57 2962 58
rect 2947 53 2948 57
rect 2952 53 2953 57
rect 2957 53 2958 57
rect 2943 52 2962 53
rect 2913 44 2915 48
rect 2919 44 2921 48
rect 2925 44 2927 48
rect 2931 44 2933 48
rect 2937 44 2939 48
rect 2943 44 2945 48
rect 2909 42 2949 44
rect 2913 38 2915 42
rect 2919 38 2921 42
rect 2925 38 2927 42
rect 2931 38 2933 42
rect 2937 38 2939 42
rect 2943 38 2945 42
rect 2909 36 2949 38
rect 2913 32 2915 36
rect 2919 32 2921 36
rect 2925 32 2927 36
rect 2931 32 2933 36
rect 2937 32 2939 36
rect 2943 32 2945 36
rect 2909 30 2949 32
rect 2913 26 2915 30
rect 2919 26 2921 30
rect 2925 26 2927 30
rect 2931 26 2933 30
rect 2937 26 2939 30
rect 2943 26 2945 30
rect 2909 24 2949 26
rect 2913 20 2915 24
rect 2919 20 2921 24
rect 2925 20 2927 24
rect 2931 20 2933 24
rect 2937 20 2939 24
rect 2943 20 2945 24
rect 2909 18 2949 20
rect 2909 14 2915 18
rect 2919 14 2921 18
rect 2925 14 2927 18
rect 2931 14 2933 18
rect 2937 14 2939 18
rect 2943 14 2945 18
rect 2909 4 2949 14
rect 2913 0 2915 4
rect 2919 0 2921 4
rect 2925 0 2927 4
rect 2931 0 2933 4
rect 2937 0 2939 4
rect 2943 0 2945 4
rect 2953 4 2962 52
rect 2986 57 3005 58
rect 2990 53 2991 57
rect 2995 53 2996 57
rect 3000 53 3001 57
rect 2986 52 3005 53
rect 2986 4 2995 52
rect 3009 48 3039 64
rect 3003 44 3005 48
rect 3009 44 3011 48
rect 3015 44 3017 48
rect 3021 44 3023 48
rect 3027 44 3029 48
rect 3033 44 3035 48
rect 2999 42 3039 44
rect 3003 38 3005 42
rect 3009 38 3011 42
rect 3015 38 3017 42
rect 3021 38 3023 42
rect 3027 38 3029 42
rect 3033 38 3035 42
rect 2999 36 3039 38
rect 3003 32 3005 36
rect 3009 32 3011 36
rect 3015 32 3017 36
rect 3021 32 3023 36
rect 3027 32 3029 36
rect 3033 32 3035 36
rect 2999 30 3039 32
rect 3003 26 3005 30
rect 3009 26 3011 30
rect 3015 26 3017 30
rect 3021 26 3023 30
rect 3027 26 3029 30
rect 3033 26 3035 30
rect 2999 24 3039 26
rect 3003 20 3005 24
rect 3009 20 3011 24
rect 3015 20 3017 24
rect 3021 20 3023 24
rect 3027 20 3029 24
rect 3033 20 3035 24
rect 2999 18 3039 20
rect 3003 14 3005 18
rect 3009 14 3011 18
rect 3015 14 3017 18
rect 3021 14 3023 18
rect 3027 14 3029 18
rect 3033 14 3039 18
rect 2999 4 3039 14
rect 3003 0 3005 4
rect 3009 0 3011 4
rect 3015 0 3017 4
rect 3021 0 3023 4
rect 3027 0 3029 4
rect 3033 0 3035 4
rect 3047 92 3049 101
rect 3053 92 3055 101
rect 3059 92 3061 101
rect 3065 92 3067 101
rect 3071 92 3073 101
rect 3077 92 3079 101
rect 3043 90 3083 92
rect 3047 86 3049 90
rect 3053 86 3055 90
rect 3059 86 3061 90
rect 3065 86 3067 90
rect 3071 86 3073 90
rect 3077 86 3079 90
rect 3043 84 3083 86
rect 3047 80 3049 84
rect 3053 80 3055 84
rect 3059 80 3061 84
rect 3065 80 3067 84
rect 3071 80 3073 84
rect 3077 80 3079 84
rect 3043 78 3083 80
rect 3047 74 3049 78
rect 3053 74 3055 78
rect 3059 74 3061 78
rect 3065 74 3067 78
rect 3071 74 3073 78
rect 3077 74 3079 78
rect 3043 72 3083 74
rect 3047 63 3049 72
rect 3053 63 3055 72
rect 3059 63 3061 72
rect 3065 63 3067 72
rect 3071 63 3073 72
rect 3077 63 3079 72
rect 3043 12 3083 63
rect 3047 8 3049 12
rect 3053 8 3055 12
rect 3059 8 3061 12
rect 3065 8 3067 12
rect 3071 8 3073 12
rect 3077 8 3079 12
rect 3043 4 3083 8
rect 3047 0 3049 4
rect 3053 0 3055 4
rect 3059 0 3061 4
rect 3065 0 3067 4
rect 3071 0 3073 4
rect 3077 0 3079 4
rect 3339 141 3379 144
rect 3343 137 3345 141
rect 3349 137 3351 141
rect 3355 137 3357 141
rect 3361 137 3363 141
rect 3367 137 3369 141
rect 3373 137 3375 141
rect 3339 101 3379 137
rect 3517 141 3557 144
rect 3521 137 3523 141
rect 3527 137 3529 141
rect 3533 137 3535 141
rect 3539 137 3541 141
rect 3545 137 3547 141
rect 3551 137 3553 141
rect 3393 131 3395 135
rect 3399 131 3401 135
rect 3405 131 3407 135
rect 3411 131 3413 135
rect 3417 131 3419 135
rect 3389 129 3423 131
rect 3387 125 3389 129
rect 3393 125 3395 129
rect 3399 125 3401 129
rect 3405 125 3407 129
rect 3411 125 3413 129
rect 3417 125 3419 129
rect 3383 123 3423 125
rect 3387 119 3389 123
rect 3393 119 3395 123
rect 3399 119 3401 123
rect 3405 119 3407 123
rect 3411 119 3413 123
rect 3417 119 3419 123
rect 3383 116 3423 119
rect 3387 112 3389 116
rect 3393 112 3395 116
rect 3399 112 3401 116
rect 3405 112 3407 116
rect 3411 112 3413 116
rect 3417 112 3419 116
rect 3383 111 3423 112
rect 3387 107 3389 111
rect 3393 107 3395 111
rect 3399 107 3401 111
rect 3405 107 3407 111
rect 3411 107 3413 111
rect 3417 107 3419 111
rect 3477 131 3479 135
rect 3483 131 3485 135
rect 3489 131 3491 135
rect 3495 131 3497 135
rect 3501 131 3503 135
rect 3473 129 3507 131
rect 3477 125 3479 129
rect 3483 125 3485 129
rect 3489 125 3491 129
rect 3495 125 3497 129
rect 3501 125 3503 129
rect 3507 125 3509 129
rect 3473 123 3513 125
rect 3477 119 3479 123
rect 3483 119 3485 123
rect 3489 119 3491 123
rect 3495 119 3497 123
rect 3501 119 3503 123
rect 3507 119 3509 123
rect 3473 116 3513 119
rect 3477 112 3479 116
rect 3483 112 3485 116
rect 3489 112 3491 116
rect 3495 112 3497 116
rect 3501 112 3503 116
rect 3507 112 3509 116
rect 3473 111 3513 112
rect 3477 107 3479 111
rect 3483 107 3485 111
rect 3489 107 3491 111
rect 3495 107 3497 111
rect 3501 107 3503 111
rect 3507 107 3509 111
rect 3343 92 3345 101
rect 3349 92 3351 101
rect 3355 92 3357 101
rect 3361 92 3363 101
rect 3367 92 3369 101
rect 3373 92 3375 101
rect 3517 101 3557 137
rect 3339 90 3379 92
rect 3343 86 3345 90
rect 3349 86 3351 90
rect 3355 86 3357 90
rect 3361 86 3363 90
rect 3367 86 3369 90
rect 3373 86 3375 90
rect 3339 84 3379 86
rect 3343 80 3345 84
rect 3349 80 3351 84
rect 3355 80 3357 84
rect 3361 80 3363 84
rect 3367 80 3369 84
rect 3373 80 3375 84
rect 3339 78 3379 80
rect 3343 74 3345 78
rect 3349 74 3351 78
rect 3355 74 3357 78
rect 3361 74 3363 78
rect 3367 74 3369 78
rect 3373 74 3375 78
rect 3339 72 3379 74
rect 3343 63 3345 72
rect 3349 63 3351 72
rect 3355 63 3357 72
rect 3361 63 3363 72
rect 3367 63 3369 72
rect 3373 63 3375 72
rect 3339 12 3379 63
rect 3343 8 3345 12
rect 3349 8 3351 12
rect 3355 8 3357 12
rect 3361 8 3363 12
rect 3367 8 3369 12
rect 3373 8 3375 12
rect 3339 4 3379 8
rect 3343 0 3345 4
rect 3349 0 3351 4
rect 3355 0 3357 4
rect 3361 0 3363 4
rect 3367 0 3369 4
rect 3373 0 3375 4
rect 3383 99 3413 100
rect 3383 95 3384 99
rect 3388 95 3390 99
rect 3394 95 3396 99
rect 3400 95 3402 99
rect 3406 95 3408 99
rect 3412 95 3413 99
rect 3383 93 3413 95
rect 3383 89 3384 93
rect 3388 89 3390 93
rect 3394 89 3396 93
rect 3400 89 3402 93
rect 3406 89 3408 93
rect 3412 89 3413 93
rect 3383 86 3413 89
rect 3383 82 3384 86
rect 3388 82 3390 86
rect 3394 82 3396 86
rect 3400 82 3402 86
rect 3406 82 3408 86
rect 3412 82 3413 86
rect 3383 80 3413 82
rect 3383 76 3384 80
rect 3388 76 3390 80
rect 3394 76 3396 80
rect 3400 76 3402 80
rect 3406 76 3408 80
rect 3412 76 3413 80
rect 3383 74 3413 76
rect 3383 70 3384 74
rect 3388 70 3390 74
rect 3394 70 3396 74
rect 3400 70 3402 74
rect 3406 70 3408 74
rect 3412 70 3413 74
rect 3383 68 3413 70
rect 3383 64 3384 68
rect 3388 64 3390 68
rect 3394 64 3396 68
rect 3400 64 3402 68
rect 3406 64 3408 68
rect 3412 64 3413 68
rect 3383 48 3413 64
rect 3483 99 3513 100
rect 3483 95 3484 99
rect 3488 95 3490 99
rect 3494 95 3496 99
rect 3500 95 3502 99
rect 3506 95 3508 99
rect 3512 95 3513 99
rect 3483 93 3513 95
rect 3483 89 3484 93
rect 3488 89 3490 93
rect 3494 89 3496 93
rect 3500 89 3502 93
rect 3506 89 3508 93
rect 3512 89 3513 93
rect 3483 86 3513 89
rect 3483 82 3484 86
rect 3488 82 3490 86
rect 3494 82 3496 86
rect 3500 82 3502 86
rect 3506 82 3508 86
rect 3512 82 3513 86
rect 3483 80 3513 82
rect 3483 76 3484 80
rect 3488 76 3490 80
rect 3494 76 3496 80
rect 3500 76 3502 80
rect 3506 76 3508 80
rect 3512 76 3513 80
rect 3483 74 3513 76
rect 3483 70 3484 74
rect 3488 70 3490 74
rect 3494 70 3496 74
rect 3500 70 3502 74
rect 3506 70 3508 74
rect 3512 70 3513 74
rect 3483 68 3513 70
rect 3483 64 3484 68
rect 3488 64 3490 68
rect 3494 64 3496 68
rect 3500 64 3502 68
rect 3506 64 3508 68
rect 3512 64 3513 68
rect 3417 57 3436 58
rect 3421 53 3422 57
rect 3426 53 3427 57
rect 3431 53 3432 57
rect 3417 52 3436 53
rect 3387 44 3389 48
rect 3393 44 3395 48
rect 3399 44 3401 48
rect 3405 44 3407 48
rect 3411 44 3413 48
rect 3417 44 3419 48
rect 3383 42 3423 44
rect 3387 38 3389 42
rect 3393 38 3395 42
rect 3399 38 3401 42
rect 3405 38 3407 42
rect 3411 38 3413 42
rect 3417 38 3419 42
rect 3383 36 3423 38
rect 3387 32 3389 36
rect 3393 32 3395 36
rect 3399 32 3401 36
rect 3405 32 3407 36
rect 3411 32 3413 36
rect 3417 32 3419 36
rect 3383 30 3423 32
rect 3387 26 3389 30
rect 3393 26 3395 30
rect 3399 26 3401 30
rect 3405 26 3407 30
rect 3411 26 3413 30
rect 3417 26 3419 30
rect 3383 24 3423 26
rect 3387 20 3389 24
rect 3393 20 3395 24
rect 3399 20 3401 24
rect 3405 20 3407 24
rect 3411 20 3413 24
rect 3417 20 3419 24
rect 3383 18 3423 20
rect 3383 14 3389 18
rect 3393 14 3395 18
rect 3399 14 3401 18
rect 3405 14 3407 18
rect 3411 14 3413 18
rect 3417 14 3419 18
rect 3383 4 3423 14
rect 3387 0 3389 4
rect 3393 0 3395 4
rect 3399 0 3401 4
rect 3405 0 3407 4
rect 3411 0 3413 4
rect 3417 0 3419 4
rect 3427 4 3436 52
rect 3460 57 3479 58
rect 3464 53 3465 57
rect 3469 53 3470 57
rect 3474 53 3475 57
rect 3460 52 3479 53
rect 3460 4 3469 52
rect 3483 48 3513 64
rect 3477 44 3479 48
rect 3483 44 3485 48
rect 3489 44 3491 48
rect 3495 44 3497 48
rect 3501 44 3503 48
rect 3507 44 3509 48
rect 3473 42 3513 44
rect 3477 38 3479 42
rect 3483 38 3485 42
rect 3489 38 3491 42
rect 3495 38 3497 42
rect 3501 38 3503 42
rect 3507 38 3509 42
rect 3473 36 3513 38
rect 3477 32 3479 36
rect 3483 32 3485 36
rect 3489 32 3491 36
rect 3495 32 3497 36
rect 3501 32 3503 36
rect 3507 32 3509 36
rect 3473 30 3513 32
rect 3477 26 3479 30
rect 3483 26 3485 30
rect 3489 26 3491 30
rect 3495 26 3497 30
rect 3501 26 3503 30
rect 3507 26 3509 30
rect 3473 24 3513 26
rect 3477 20 3479 24
rect 3483 20 3485 24
rect 3489 20 3491 24
rect 3495 20 3497 24
rect 3501 20 3503 24
rect 3507 20 3509 24
rect 3473 18 3513 20
rect 3477 14 3479 18
rect 3483 14 3485 18
rect 3489 14 3491 18
rect 3495 14 3497 18
rect 3501 14 3503 18
rect 3507 14 3513 18
rect 3473 4 3513 14
rect 3477 0 3479 4
rect 3483 0 3485 4
rect 3489 0 3491 4
rect 3495 0 3497 4
rect 3501 0 3503 4
rect 3507 0 3509 4
rect 3521 92 3523 101
rect 3527 92 3529 101
rect 3533 92 3535 101
rect 3539 92 3541 101
rect 3545 92 3547 101
rect 3551 92 3553 101
rect 3517 90 3557 92
rect 3521 86 3523 90
rect 3527 86 3529 90
rect 3533 86 3535 90
rect 3539 86 3541 90
rect 3545 86 3547 90
rect 3551 86 3553 90
rect 3517 84 3557 86
rect 3521 80 3523 84
rect 3527 80 3529 84
rect 3533 80 3535 84
rect 3539 80 3541 84
rect 3545 80 3547 84
rect 3551 80 3553 84
rect 3517 78 3557 80
rect 3521 74 3523 78
rect 3527 74 3529 78
rect 3533 74 3535 78
rect 3539 74 3541 78
rect 3545 74 3547 78
rect 3551 74 3553 78
rect 3517 72 3557 74
rect 3521 63 3523 72
rect 3527 63 3529 72
rect 3533 63 3535 72
rect 3539 63 3541 72
rect 3545 63 3547 72
rect 3551 63 3553 72
rect 3517 12 3557 63
rect 3521 8 3523 12
rect 3527 8 3529 12
rect 3533 8 3535 12
rect 3539 8 3541 12
rect 3545 8 3547 12
rect 3551 8 3553 12
rect 3517 4 3557 8
rect 3521 0 3523 4
rect 3527 0 3529 4
rect 3533 0 3535 4
rect 3539 0 3541 4
rect 3545 0 3547 4
rect 3551 0 3553 4
rect 3813 141 3853 144
rect 3817 137 3819 141
rect 3823 137 3825 141
rect 3829 137 3831 141
rect 3835 137 3837 141
rect 3841 137 3843 141
rect 3847 137 3849 141
rect 3813 101 3853 137
rect 3991 141 4031 144
rect 3995 137 3997 141
rect 4001 137 4003 141
rect 4007 137 4009 141
rect 4013 137 4015 141
rect 4019 137 4021 141
rect 4025 137 4027 141
rect 3867 131 3869 135
rect 3873 131 3875 135
rect 3879 131 3881 135
rect 3885 131 3887 135
rect 3891 131 3893 135
rect 3863 129 3897 131
rect 3861 125 3863 129
rect 3867 125 3869 129
rect 3873 125 3875 129
rect 3879 125 3881 129
rect 3885 125 3887 129
rect 3891 125 3893 129
rect 3857 123 3897 125
rect 3861 119 3863 123
rect 3867 119 3869 123
rect 3873 119 3875 123
rect 3879 119 3881 123
rect 3885 119 3887 123
rect 3891 119 3893 123
rect 3857 116 3897 119
rect 3861 112 3863 116
rect 3867 112 3869 116
rect 3873 112 3875 116
rect 3879 112 3881 116
rect 3885 112 3887 116
rect 3891 112 3893 116
rect 3857 111 3897 112
rect 3861 107 3863 111
rect 3867 107 3869 111
rect 3873 107 3875 111
rect 3879 107 3881 111
rect 3885 107 3887 111
rect 3891 107 3893 111
rect 3951 131 3953 135
rect 3957 131 3959 135
rect 3963 131 3965 135
rect 3969 131 3971 135
rect 3975 131 3977 135
rect 3947 129 3981 131
rect 3951 125 3953 129
rect 3957 125 3959 129
rect 3963 125 3965 129
rect 3969 125 3971 129
rect 3975 125 3977 129
rect 3981 125 3983 129
rect 3947 123 3987 125
rect 3951 119 3953 123
rect 3957 119 3959 123
rect 3963 119 3965 123
rect 3969 119 3971 123
rect 3975 119 3977 123
rect 3981 119 3983 123
rect 3947 116 3987 119
rect 3951 112 3953 116
rect 3957 112 3959 116
rect 3963 112 3965 116
rect 3969 112 3971 116
rect 3975 112 3977 116
rect 3981 112 3983 116
rect 3947 111 3987 112
rect 3951 107 3953 111
rect 3957 107 3959 111
rect 3963 107 3965 111
rect 3969 107 3971 111
rect 3975 107 3977 111
rect 3981 107 3983 111
rect 3817 92 3819 101
rect 3823 92 3825 101
rect 3829 92 3831 101
rect 3835 92 3837 101
rect 3841 92 3843 101
rect 3847 92 3849 101
rect 3991 101 4031 137
rect 3813 90 3853 92
rect 3817 86 3819 90
rect 3823 86 3825 90
rect 3829 86 3831 90
rect 3835 86 3837 90
rect 3841 86 3843 90
rect 3847 86 3849 90
rect 3813 84 3853 86
rect 3817 80 3819 84
rect 3823 80 3825 84
rect 3829 80 3831 84
rect 3835 80 3837 84
rect 3841 80 3843 84
rect 3847 80 3849 84
rect 3813 78 3853 80
rect 3817 74 3819 78
rect 3823 74 3825 78
rect 3829 74 3831 78
rect 3835 74 3837 78
rect 3841 74 3843 78
rect 3847 74 3849 78
rect 3813 72 3853 74
rect 3817 63 3819 72
rect 3823 63 3825 72
rect 3829 63 3831 72
rect 3835 63 3837 72
rect 3841 63 3843 72
rect 3847 63 3849 72
rect 3813 12 3853 63
rect 3817 8 3819 12
rect 3823 8 3825 12
rect 3829 8 3831 12
rect 3835 8 3837 12
rect 3841 8 3843 12
rect 3847 8 3849 12
rect 3813 4 3853 8
rect 3817 0 3819 4
rect 3823 0 3825 4
rect 3829 0 3831 4
rect 3835 0 3837 4
rect 3841 0 3843 4
rect 3847 0 3849 4
rect 3857 99 3887 100
rect 3857 95 3858 99
rect 3862 95 3864 99
rect 3868 95 3870 99
rect 3874 95 3876 99
rect 3880 95 3882 99
rect 3886 95 3887 99
rect 3857 93 3887 95
rect 3857 89 3858 93
rect 3862 89 3864 93
rect 3868 89 3870 93
rect 3874 89 3876 93
rect 3880 89 3882 93
rect 3886 89 3887 93
rect 3857 86 3887 89
rect 3857 82 3858 86
rect 3862 82 3864 86
rect 3868 82 3870 86
rect 3874 82 3876 86
rect 3880 82 3882 86
rect 3886 82 3887 86
rect 3857 80 3887 82
rect 3857 76 3858 80
rect 3862 76 3864 80
rect 3868 76 3870 80
rect 3874 76 3876 80
rect 3880 76 3882 80
rect 3886 76 3887 80
rect 3857 74 3887 76
rect 3857 70 3858 74
rect 3862 70 3864 74
rect 3868 70 3870 74
rect 3874 70 3876 74
rect 3880 70 3882 74
rect 3886 70 3887 74
rect 3857 68 3887 70
rect 3857 64 3858 68
rect 3862 64 3864 68
rect 3868 64 3870 68
rect 3874 64 3876 68
rect 3880 64 3882 68
rect 3886 64 3887 68
rect 3857 48 3887 64
rect 3957 99 3987 100
rect 3957 95 3958 99
rect 3962 95 3964 99
rect 3968 95 3970 99
rect 3974 95 3976 99
rect 3980 95 3982 99
rect 3986 95 3987 99
rect 3957 93 3987 95
rect 3957 89 3958 93
rect 3962 89 3964 93
rect 3968 89 3970 93
rect 3974 89 3976 93
rect 3980 89 3982 93
rect 3986 89 3987 93
rect 3957 86 3987 89
rect 3957 82 3958 86
rect 3962 82 3964 86
rect 3968 82 3970 86
rect 3974 82 3976 86
rect 3980 82 3982 86
rect 3986 82 3987 86
rect 3957 80 3987 82
rect 3957 76 3958 80
rect 3962 76 3964 80
rect 3968 76 3970 80
rect 3974 76 3976 80
rect 3980 76 3982 80
rect 3986 76 3987 80
rect 3957 74 3987 76
rect 3957 70 3958 74
rect 3962 70 3964 74
rect 3968 70 3970 74
rect 3974 70 3976 74
rect 3980 70 3982 74
rect 3986 70 3987 74
rect 3957 68 3987 70
rect 3957 64 3958 68
rect 3962 64 3964 68
rect 3968 64 3970 68
rect 3974 64 3976 68
rect 3980 64 3982 68
rect 3986 64 3987 68
rect 3891 57 3910 58
rect 3895 53 3896 57
rect 3900 53 3901 57
rect 3905 53 3906 57
rect 3891 52 3910 53
rect 3861 44 3863 48
rect 3867 44 3869 48
rect 3873 44 3875 48
rect 3879 44 3881 48
rect 3885 44 3887 48
rect 3891 44 3893 48
rect 3857 42 3897 44
rect 3861 38 3863 42
rect 3867 38 3869 42
rect 3873 38 3875 42
rect 3879 38 3881 42
rect 3885 38 3887 42
rect 3891 38 3893 42
rect 3857 36 3897 38
rect 3861 32 3863 36
rect 3867 32 3869 36
rect 3873 32 3875 36
rect 3879 32 3881 36
rect 3885 32 3887 36
rect 3891 32 3893 36
rect 3857 30 3897 32
rect 3861 26 3863 30
rect 3867 26 3869 30
rect 3873 26 3875 30
rect 3879 26 3881 30
rect 3885 26 3887 30
rect 3891 26 3893 30
rect 3857 24 3897 26
rect 3861 20 3863 24
rect 3867 20 3869 24
rect 3873 20 3875 24
rect 3879 20 3881 24
rect 3885 20 3887 24
rect 3891 20 3893 24
rect 3857 18 3897 20
rect 3857 14 3863 18
rect 3867 14 3869 18
rect 3873 14 3875 18
rect 3879 14 3881 18
rect 3885 14 3887 18
rect 3891 14 3893 18
rect 3857 4 3897 14
rect 3861 0 3863 4
rect 3867 0 3869 4
rect 3873 0 3875 4
rect 3879 0 3881 4
rect 3885 0 3887 4
rect 3891 0 3893 4
rect 3901 4 3910 52
rect 3934 57 3953 58
rect 3938 53 3939 57
rect 3943 53 3944 57
rect 3948 53 3949 57
rect 3934 52 3953 53
rect 3934 4 3943 52
rect 3957 48 3987 64
rect 3951 44 3953 48
rect 3957 44 3959 48
rect 3963 44 3965 48
rect 3969 44 3971 48
rect 3975 44 3977 48
rect 3981 44 3983 48
rect 3947 42 3987 44
rect 3951 38 3953 42
rect 3957 38 3959 42
rect 3963 38 3965 42
rect 3969 38 3971 42
rect 3975 38 3977 42
rect 3981 38 3983 42
rect 3947 36 3987 38
rect 3951 32 3953 36
rect 3957 32 3959 36
rect 3963 32 3965 36
rect 3969 32 3971 36
rect 3975 32 3977 36
rect 3981 32 3983 36
rect 3947 30 3987 32
rect 3951 26 3953 30
rect 3957 26 3959 30
rect 3963 26 3965 30
rect 3969 26 3971 30
rect 3975 26 3977 30
rect 3981 26 3983 30
rect 3947 24 3987 26
rect 3951 20 3953 24
rect 3957 20 3959 24
rect 3963 20 3965 24
rect 3969 20 3971 24
rect 3975 20 3977 24
rect 3981 20 3983 24
rect 3947 18 3987 20
rect 3951 14 3953 18
rect 3957 14 3959 18
rect 3963 14 3965 18
rect 3969 14 3971 18
rect 3975 14 3977 18
rect 3981 14 3987 18
rect 3947 4 3987 14
rect 3951 0 3953 4
rect 3957 0 3959 4
rect 3963 0 3965 4
rect 3969 0 3971 4
rect 3975 0 3977 4
rect 3981 0 3983 4
rect 3995 92 3997 101
rect 4001 92 4003 101
rect 4007 92 4009 101
rect 4013 92 4015 101
rect 4019 92 4021 101
rect 4025 92 4027 101
rect 3991 90 4031 92
rect 3995 86 3997 90
rect 4001 86 4003 90
rect 4007 86 4009 90
rect 4013 86 4015 90
rect 4019 86 4021 90
rect 4025 86 4027 90
rect 3991 84 4031 86
rect 3995 80 3997 84
rect 4001 80 4003 84
rect 4007 80 4009 84
rect 4013 80 4015 84
rect 4019 80 4021 84
rect 4025 80 4027 84
rect 3991 78 4031 80
rect 3995 74 3997 78
rect 4001 74 4003 78
rect 4007 74 4009 78
rect 4013 74 4015 78
rect 4019 74 4021 78
rect 4025 74 4027 78
rect 3991 72 4031 74
rect 3995 63 3997 72
rect 4001 63 4003 72
rect 4007 63 4009 72
rect 4013 63 4015 72
rect 4019 63 4021 72
rect 4025 63 4027 72
rect 3991 12 4031 63
rect 3995 8 3997 12
rect 4001 8 4003 12
rect 4007 8 4009 12
rect 4013 8 4015 12
rect 4019 8 4021 12
rect 4025 8 4027 12
rect 3991 4 4031 8
rect 3995 0 3997 4
rect 4001 0 4003 4
rect 4007 0 4009 4
rect 4013 0 4015 4
rect 4019 0 4021 4
rect 4025 0 4027 4
rect 4287 141 4327 144
rect 4291 137 4293 141
rect 4297 137 4299 141
rect 4303 137 4305 141
rect 4309 137 4311 141
rect 4315 137 4317 141
rect 4321 137 4323 141
rect 4287 101 4327 137
rect 4465 141 4505 144
rect 4469 137 4471 141
rect 4475 137 4477 141
rect 4481 137 4483 141
rect 4487 137 4489 141
rect 4493 137 4495 141
rect 4499 137 4501 141
rect 4341 131 4343 135
rect 4347 131 4349 135
rect 4353 131 4355 135
rect 4359 131 4361 135
rect 4365 131 4367 135
rect 4337 129 4371 131
rect 4335 125 4337 129
rect 4341 125 4343 129
rect 4347 125 4349 129
rect 4353 125 4355 129
rect 4359 125 4361 129
rect 4365 125 4367 129
rect 4331 123 4371 125
rect 4335 119 4337 123
rect 4341 119 4343 123
rect 4347 119 4349 123
rect 4353 119 4355 123
rect 4359 119 4361 123
rect 4365 119 4367 123
rect 4331 116 4371 119
rect 4335 112 4337 116
rect 4341 112 4343 116
rect 4347 112 4349 116
rect 4353 112 4355 116
rect 4359 112 4361 116
rect 4365 112 4367 116
rect 4331 111 4371 112
rect 4335 107 4337 111
rect 4341 107 4343 111
rect 4347 107 4349 111
rect 4353 107 4355 111
rect 4359 107 4361 111
rect 4365 107 4367 111
rect 4425 131 4427 135
rect 4431 131 4433 135
rect 4437 131 4439 135
rect 4443 131 4445 135
rect 4449 131 4451 135
rect 4421 129 4455 131
rect 4425 125 4427 129
rect 4431 125 4433 129
rect 4437 125 4439 129
rect 4443 125 4445 129
rect 4449 125 4451 129
rect 4455 125 4457 129
rect 4421 123 4461 125
rect 4425 119 4427 123
rect 4431 119 4433 123
rect 4437 119 4439 123
rect 4443 119 4445 123
rect 4449 119 4451 123
rect 4455 119 4457 123
rect 4421 116 4461 119
rect 4425 112 4427 116
rect 4431 112 4433 116
rect 4437 112 4439 116
rect 4443 112 4445 116
rect 4449 112 4451 116
rect 4455 112 4457 116
rect 4421 111 4461 112
rect 4425 107 4427 111
rect 4431 107 4433 111
rect 4437 107 4439 111
rect 4443 107 4445 111
rect 4449 107 4451 111
rect 4455 107 4457 111
rect 4291 92 4293 101
rect 4297 92 4299 101
rect 4303 92 4305 101
rect 4309 92 4311 101
rect 4315 92 4317 101
rect 4321 92 4323 101
rect 4465 101 4505 137
rect 4287 90 4327 92
rect 4291 86 4293 90
rect 4297 86 4299 90
rect 4303 86 4305 90
rect 4309 86 4311 90
rect 4315 86 4317 90
rect 4321 86 4323 90
rect 4287 84 4327 86
rect 4291 80 4293 84
rect 4297 80 4299 84
rect 4303 80 4305 84
rect 4309 80 4311 84
rect 4315 80 4317 84
rect 4321 80 4323 84
rect 4287 78 4327 80
rect 4291 74 4293 78
rect 4297 74 4299 78
rect 4303 74 4305 78
rect 4309 74 4311 78
rect 4315 74 4317 78
rect 4321 74 4323 78
rect 4287 72 4327 74
rect 4291 63 4293 72
rect 4297 63 4299 72
rect 4303 63 4305 72
rect 4309 63 4311 72
rect 4315 63 4317 72
rect 4321 63 4323 72
rect 4287 12 4327 63
rect 4291 8 4293 12
rect 4297 8 4299 12
rect 4303 8 4305 12
rect 4309 8 4311 12
rect 4315 8 4317 12
rect 4321 8 4323 12
rect 4287 4 4327 8
rect 4291 0 4293 4
rect 4297 0 4299 4
rect 4303 0 4305 4
rect 4309 0 4311 4
rect 4315 0 4317 4
rect 4321 0 4323 4
rect 4331 99 4361 100
rect 4331 95 4332 99
rect 4336 95 4338 99
rect 4342 95 4344 99
rect 4348 95 4350 99
rect 4354 95 4356 99
rect 4360 95 4361 99
rect 4331 93 4361 95
rect 4331 89 4332 93
rect 4336 89 4338 93
rect 4342 89 4344 93
rect 4348 89 4350 93
rect 4354 89 4356 93
rect 4360 89 4361 93
rect 4331 86 4361 89
rect 4331 82 4332 86
rect 4336 82 4338 86
rect 4342 82 4344 86
rect 4348 82 4350 86
rect 4354 82 4356 86
rect 4360 82 4361 86
rect 4331 80 4361 82
rect 4331 76 4332 80
rect 4336 76 4338 80
rect 4342 76 4344 80
rect 4348 76 4350 80
rect 4354 76 4356 80
rect 4360 76 4361 80
rect 4331 74 4361 76
rect 4331 70 4332 74
rect 4336 70 4338 74
rect 4342 70 4344 74
rect 4348 70 4350 74
rect 4354 70 4356 74
rect 4360 70 4361 74
rect 4331 68 4361 70
rect 4331 64 4332 68
rect 4336 64 4338 68
rect 4342 64 4344 68
rect 4348 64 4350 68
rect 4354 64 4356 68
rect 4360 64 4361 68
rect 4331 48 4361 64
rect 4431 99 4461 100
rect 4431 95 4432 99
rect 4436 95 4438 99
rect 4442 95 4444 99
rect 4448 95 4450 99
rect 4454 95 4456 99
rect 4460 95 4461 99
rect 4431 93 4461 95
rect 4431 89 4432 93
rect 4436 89 4438 93
rect 4442 89 4444 93
rect 4448 89 4450 93
rect 4454 89 4456 93
rect 4460 89 4461 93
rect 4431 86 4461 89
rect 4431 82 4432 86
rect 4436 82 4438 86
rect 4442 82 4444 86
rect 4448 82 4450 86
rect 4454 82 4456 86
rect 4460 82 4461 86
rect 4431 80 4461 82
rect 4431 76 4432 80
rect 4436 76 4438 80
rect 4442 76 4444 80
rect 4448 76 4450 80
rect 4454 76 4456 80
rect 4460 76 4461 80
rect 4431 74 4461 76
rect 4431 70 4432 74
rect 4436 70 4438 74
rect 4442 70 4444 74
rect 4448 70 4450 74
rect 4454 70 4456 74
rect 4460 70 4461 74
rect 4431 68 4461 70
rect 4431 64 4432 68
rect 4436 64 4438 68
rect 4442 64 4444 68
rect 4448 64 4450 68
rect 4454 64 4456 68
rect 4460 64 4461 68
rect 4365 57 4384 58
rect 4369 53 4370 57
rect 4374 53 4375 57
rect 4379 53 4380 57
rect 4365 52 4384 53
rect 4335 44 4337 48
rect 4341 44 4343 48
rect 4347 44 4349 48
rect 4353 44 4355 48
rect 4359 44 4361 48
rect 4365 44 4367 48
rect 4331 42 4371 44
rect 4335 38 4337 42
rect 4341 38 4343 42
rect 4347 38 4349 42
rect 4353 38 4355 42
rect 4359 38 4361 42
rect 4365 38 4367 42
rect 4331 36 4371 38
rect 4335 32 4337 36
rect 4341 32 4343 36
rect 4347 32 4349 36
rect 4353 32 4355 36
rect 4359 32 4361 36
rect 4365 32 4367 36
rect 4331 30 4371 32
rect 4335 26 4337 30
rect 4341 26 4343 30
rect 4347 26 4349 30
rect 4353 26 4355 30
rect 4359 26 4361 30
rect 4365 26 4367 30
rect 4331 24 4371 26
rect 4335 20 4337 24
rect 4341 20 4343 24
rect 4347 20 4349 24
rect 4353 20 4355 24
rect 4359 20 4361 24
rect 4365 20 4367 24
rect 4331 18 4371 20
rect 4331 14 4337 18
rect 4341 14 4343 18
rect 4347 14 4349 18
rect 4353 14 4355 18
rect 4359 14 4361 18
rect 4365 14 4367 18
rect 4331 4 4371 14
rect 4335 0 4337 4
rect 4341 0 4343 4
rect 4347 0 4349 4
rect 4353 0 4355 4
rect 4359 0 4361 4
rect 4365 0 4367 4
rect 4375 4 4384 52
rect 4408 57 4427 58
rect 4412 53 4413 57
rect 4417 53 4418 57
rect 4422 53 4423 57
rect 4408 52 4427 53
rect 4408 4 4417 52
rect 4431 48 4461 64
rect 4469 92 4471 101
rect 4475 92 4477 101
rect 4481 92 4483 101
rect 4487 92 4489 101
rect 4493 92 4495 101
rect 4499 92 4501 101
rect 4465 90 4505 92
rect 4469 86 4471 90
rect 4475 86 4477 90
rect 4481 86 4483 90
rect 4487 86 4489 90
rect 4493 86 4495 90
rect 4499 86 4501 90
rect 4465 84 4505 86
rect 4469 80 4471 84
rect 4475 80 4477 84
rect 4481 80 4483 84
rect 4487 80 4489 84
rect 4493 80 4495 84
rect 4499 80 4501 84
rect 4465 78 4505 80
rect 4469 74 4471 78
rect 4475 74 4477 78
rect 4481 74 4483 78
rect 4487 74 4489 78
rect 4493 74 4495 78
rect 4499 74 4501 78
rect 4465 72 4505 74
rect 4469 63 4471 72
rect 4475 63 4477 72
rect 4481 63 4483 72
rect 4487 63 4489 72
rect 4493 63 4495 72
rect 4499 63 4501 72
rect 4465 62 4505 63
rect 4425 44 4427 48
rect 4431 44 4433 48
rect 4437 44 4439 48
rect 4443 44 4445 48
rect 4449 44 4451 48
rect 4455 44 4457 48
rect 4421 42 4461 44
rect 4425 38 4427 42
rect 4431 38 4433 42
rect 4437 38 4439 42
rect 4443 38 4445 42
rect 4449 38 4451 42
rect 4455 38 4457 42
rect 4421 36 4461 38
rect 4425 32 4427 36
rect 4431 32 4433 36
rect 4437 32 4439 36
rect 4443 32 4445 36
rect 4449 32 4451 36
rect 4455 32 4457 36
rect 4421 30 4461 32
rect 4425 26 4427 30
rect 4431 26 4433 30
rect 4437 26 4439 30
rect 4443 26 4445 30
rect 4449 26 4451 30
rect 4455 26 4457 30
rect 4421 24 4461 26
rect 4425 20 4427 24
rect 4431 20 4433 24
rect 4437 20 4439 24
rect 4443 20 4445 24
rect 4449 20 4451 24
rect 4455 20 4457 24
rect 4421 18 4461 20
rect 4425 14 4427 18
rect 4431 14 4433 18
rect 4437 14 4439 18
rect 4443 14 4445 18
rect 4449 14 4451 18
rect 4455 14 4457 18
rect 4421 4 4461 14
rect 4425 0 4427 4
rect 4431 0 4433 4
rect 4437 0 4439 4
rect 4443 0 4445 4
rect 4449 0 4451 4
rect 4455 0 4457 4
<< m2contact >>
rect 4654 490 4668 499
rect 4643 176 4647 180
rect 4643 168 4647 172
rect 4675 176 4679 180
rect 4675 168 4679 172
rect 4643 160 4647 164
rect 4675 160 4679 164
rect 4651 156 4655 160
rect 4659 156 4663 160
rect 4667 156 4671 160
rect 4699 176 4703 180
rect 4699 168 4703 172
rect 4731 176 4735 180
rect 4731 168 4735 172
rect 4699 160 4703 164
rect 4731 160 4735 164
rect 4707 156 4711 160
rect 4715 156 4719 160
rect 4723 156 4727 160
rect 545 131 549 135
rect 551 131 555 135
rect 557 131 561 135
rect 563 131 567 135
rect 569 131 573 135
rect 575 131 579 135
rect 539 119 543 123
rect 545 119 549 123
rect 551 119 555 123
rect 557 119 561 123
rect 563 119 567 123
rect 569 119 573 123
rect 575 119 579 123
rect 539 107 543 111
rect 545 107 549 111
rect 551 107 555 111
rect 557 107 561 111
rect 563 107 567 111
rect 569 107 573 111
rect 575 107 579 111
rect 629 131 633 135
rect 635 131 639 135
rect 641 131 645 135
rect 647 131 651 135
rect 653 131 657 135
rect 659 131 663 135
rect 629 119 633 123
rect 635 119 639 123
rect 641 119 645 123
rect 647 119 651 123
rect 653 119 657 123
rect 659 119 663 123
rect 665 119 669 123
rect 629 107 633 111
rect 635 107 639 111
rect 641 107 645 111
rect 647 107 651 111
rect 653 107 657 111
rect 659 107 663 111
rect 665 107 669 111
rect 495 92 499 101
rect 501 92 505 101
rect 507 92 511 101
rect 513 92 517 101
rect 519 92 523 101
rect 525 92 529 101
rect 531 92 535 101
rect 495 86 499 90
rect 501 86 505 90
rect 507 86 511 90
rect 513 86 517 90
rect 519 86 523 90
rect 525 86 529 90
rect 531 86 535 90
rect 495 80 499 84
rect 501 80 505 84
rect 507 80 511 84
rect 513 80 517 84
rect 519 80 523 84
rect 525 80 529 84
rect 531 80 535 84
rect 495 74 499 78
rect 501 74 505 78
rect 507 74 511 78
rect 513 74 517 78
rect 519 74 523 78
rect 525 74 529 78
rect 531 74 535 78
rect 495 63 499 72
rect 501 63 505 72
rect 507 63 511 72
rect 513 63 517 72
rect 519 63 523 72
rect 525 63 529 72
rect 531 63 535 72
rect 578 53 582 57
rect 588 53 592 57
rect 539 43 543 47
rect 545 43 549 47
rect 551 43 555 47
rect 557 43 561 47
rect 563 43 567 47
rect 569 43 573 47
rect 575 43 579 47
rect 539 32 543 36
rect 545 32 549 36
rect 551 32 555 36
rect 557 32 561 36
rect 563 32 567 36
rect 569 32 573 36
rect 575 32 579 36
rect 539 26 543 30
rect 545 26 549 30
rect 551 26 555 30
rect 557 26 561 30
rect 563 26 567 30
rect 569 26 573 30
rect 575 26 579 30
rect 539 14 543 18
rect 545 14 549 18
rect 551 14 555 18
rect 557 14 561 18
rect 563 14 567 18
rect 569 14 573 18
rect 575 14 579 18
rect 539 0 543 4
rect 545 0 549 4
rect 551 0 555 4
rect 557 0 561 4
rect 563 0 567 4
rect 569 0 573 4
rect 575 0 579 4
rect 583 0 592 4
rect 616 53 620 57
rect 626 53 630 57
rect 616 0 625 4
rect 629 43 633 47
rect 635 43 639 47
rect 641 43 645 47
rect 647 43 651 47
rect 653 43 657 47
rect 659 43 663 47
rect 665 43 669 47
rect 629 32 633 36
rect 635 32 639 36
rect 641 32 645 36
rect 647 32 651 36
rect 653 32 657 36
rect 659 32 663 36
rect 665 32 669 36
rect 629 26 633 30
rect 635 26 639 30
rect 641 26 645 30
rect 647 26 651 30
rect 653 26 657 30
rect 659 26 663 30
rect 665 26 669 30
rect 629 14 633 18
rect 635 14 639 18
rect 641 14 645 18
rect 647 14 651 18
rect 653 14 657 18
rect 659 14 663 18
rect 629 0 633 4
rect 635 0 639 4
rect 641 0 645 4
rect 647 0 651 4
rect 653 0 657 4
rect 659 0 663 4
rect 665 0 669 4
rect 673 92 677 101
rect 679 92 683 101
rect 685 92 689 101
rect 691 92 695 101
rect 697 92 701 101
rect 703 92 707 101
rect 709 92 713 101
rect 673 86 677 90
rect 679 86 683 90
rect 685 86 689 90
rect 691 86 695 90
rect 697 86 701 90
rect 703 86 707 90
rect 709 86 713 90
rect 673 80 677 84
rect 679 80 683 84
rect 685 80 689 84
rect 691 80 695 84
rect 697 80 701 84
rect 703 80 707 84
rect 709 80 713 84
rect 673 74 677 78
rect 679 74 683 78
rect 685 74 689 78
rect 691 74 695 78
rect 697 74 701 78
rect 703 74 707 78
rect 709 74 713 78
rect 673 63 677 72
rect 679 63 683 72
rect 685 63 689 72
rect 691 63 695 72
rect 697 63 701 72
rect 703 63 707 72
rect 709 63 713 72
rect 673 0 677 4
rect 679 0 683 4
rect 685 0 689 4
rect 691 0 695 4
rect 697 0 701 4
rect 703 0 707 4
rect 709 0 713 4
rect 1019 131 1023 135
rect 1025 131 1029 135
rect 1031 131 1035 135
rect 1037 131 1041 135
rect 1043 131 1047 135
rect 1049 131 1053 135
rect 1013 119 1017 123
rect 1019 119 1023 123
rect 1025 119 1029 123
rect 1031 119 1035 123
rect 1037 119 1041 123
rect 1043 119 1047 123
rect 1049 119 1053 123
rect 1013 107 1017 111
rect 1019 107 1023 111
rect 1025 107 1029 111
rect 1031 107 1035 111
rect 1037 107 1041 111
rect 1043 107 1047 111
rect 1049 107 1053 111
rect 1103 131 1107 135
rect 1109 131 1113 135
rect 1115 131 1119 135
rect 1121 131 1125 135
rect 1127 131 1131 135
rect 1133 131 1137 135
rect 1103 119 1107 123
rect 1109 119 1113 123
rect 1115 119 1119 123
rect 1121 119 1125 123
rect 1127 119 1131 123
rect 1133 119 1137 123
rect 1139 119 1143 123
rect 1103 107 1107 111
rect 1109 107 1113 111
rect 1115 107 1119 111
rect 1121 107 1125 111
rect 1127 107 1131 111
rect 1133 107 1137 111
rect 1139 107 1143 111
rect 969 92 973 101
rect 975 92 979 101
rect 981 92 985 101
rect 987 92 991 101
rect 993 92 997 101
rect 999 92 1003 101
rect 1005 92 1009 101
rect 969 86 973 90
rect 975 86 979 90
rect 981 86 985 90
rect 987 86 991 90
rect 993 86 997 90
rect 999 86 1003 90
rect 1005 86 1009 90
rect 969 80 973 84
rect 975 80 979 84
rect 981 80 985 84
rect 987 80 991 84
rect 993 80 997 84
rect 999 80 1003 84
rect 1005 80 1009 84
rect 969 74 973 78
rect 975 74 979 78
rect 981 74 985 78
rect 987 74 991 78
rect 993 74 997 78
rect 999 74 1003 78
rect 1005 74 1009 78
rect 969 63 973 72
rect 975 63 979 72
rect 981 63 985 72
rect 987 63 991 72
rect 993 63 997 72
rect 999 63 1003 72
rect 1005 63 1009 72
rect 969 0 973 4
rect 975 0 979 4
rect 981 0 985 4
rect 987 0 991 4
rect 993 0 997 4
rect 999 0 1003 4
rect 1005 0 1009 4
rect 1052 53 1056 57
rect 1062 53 1066 57
rect 1013 44 1017 48
rect 1019 44 1023 48
rect 1025 44 1029 48
rect 1031 44 1035 48
rect 1037 44 1041 48
rect 1043 44 1047 48
rect 1049 44 1053 48
rect 1013 32 1017 36
rect 1019 32 1023 36
rect 1025 32 1029 36
rect 1031 32 1035 36
rect 1037 32 1041 36
rect 1043 32 1047 36
rect 1049 32 1053 36
rect 1013 26 1017 30
rect 1019 26 1023 30
rect 1025 26 1029 30
rect 1031 26 1035 30
rect 1037 26 1041 30
rect 1043 26 1047 30
rect 1049 26 1053 30
rect 1019 14 1023 18
rect 1025 14 1029 18
rect 1031 14 1035 18
rect 1037 14 1041 18
rect 1043 14 1047 18
rect 1049 14 1053 18
rect 1013 0 1017 4
rect 1019 0 1023 4
rect 1025 0 1029 4
rect 1031 0 1035 4
rect 1037 0 1041 4
rect 1043 0 1047 4
rect 1049 0 1053 4
rect 1057 0 1066 4
rect 1090 53 1094 57
rect 1100 53 1104 57
rect 1090 0 1099 4
rect 1103 44 1107 48
rect 1109 44 1113 48
rect 1115 44 1119 48
rect 1121 44 1125 48
rect 1127 44 1131 48
rect 1133 44 1137 48
rect 1139 44 1143 48
rect 1103 32 1107 36
rect 1109 32 1113 36
rect 1115 32 1119 36
rect 1121 32 1125 36
rect 1127 32 1131 36
rect 1133 32 1137 36
rect 1139 32 1143 36
rect 1103 26 1107 30
rect 1109 26 1113 30
rect 1115 26 1119 30
rect 1121 26 1125 30
rect 1127 26 1131 30
rect 1133 26 1137 30
rect 1139 26 1143 30
rect 1103 14 1107 18
rect 1109 14 1113 18
rect 1115 14 1119 18
rect 1121 14 1125 18
rect 1127 14 1131 18
rect 1133 14 1137 18
rect 1103 0 1107 4
rect 1109 0 1113 4
rect 1115 0 1119 4
rect 1121 0 1125 4
rect 1127 0 1131 4
rect 1133 0 1137 4
rect 1139 0 1143 4
rect 1147 92 1151 101
rect 1153 92 1157 101
rect 1159 92 1163 101
rect 1165 92 1169 101
rect 1171 92 1175 101
rect 1177 92 1181 101
rect 1183 92 1187 101
rect 1147 86 1151 90
rect 1153 86 1157 90
rect 1159 86 1163 90
rect 1165 86 1169 90
rect 1171 86 1175 90
rect 1177 86 1181 90
rect 1183 86 1187 90
rect 1147 80 1151 84
rect 1153 80 1157 84
rect 1159 80 1163 84
rect 1165 80 1169 84
rect 1171 80 1175 84
rect 1177 80 1181 84
rect 1183 80 1187 84
rect 1147 74 1151 78
rect 1153 74 1157 78
rect 1159 74 1163 78
rect 1165 74 1169 78
rect 1171 74 1175 78
rect 1177 74 1181 78
rect 1183 74 1187 78
rect 1147 63 1151 72
rect 1153 63 1157 72
rect 1159 63 1163 72
rect 1165 63 1169 72
rect 1171 63 1175 72
rect 1177 63 1181 72
rect 1183 63 1187 72
rect 1147 0 1151 4
rect 1153 0 1157 4
rect 1159 0 1163 4
rect 1165 0 1169 4
rect 1171 0 1175 4
rect 1177 0 1181 4
rect 1183 0 1187 4
rect 1493 131 1497 135
rect 1499 131 1503 135
rect 1505 131 1509 135
rect 1511 131 1515 135
rect 1517 131 1521 135
rect 1523 131 1527 135
rect 1487 119 1491 123
rect 1493 119 1497 123
rect 1499 119 1503 123
rect 1505 119 1509 123
rect 1511 119 1515 123
rect 1517 119 1521 123
rect 1523 119 1527 123
rect 1487 107 1491 111
rect 1493 107 1497 111
rect 1499 107 1503 111
rect 1505 107 1509 111
rect 1511 107 1515 111
rect 1517 107 1521 111
rect 1523 107 1527 111
rect 1577 131 1581 135
rect 1583 131 1587 135
rect 1589 131 1593 135
rect 1595 131 1599 135
rect 1601 131 1605 135
rect 1607 131 1611 135
rect 1577 119 1581 123
rect 1583 119 1587 123
rect 1589 119 1593 123
rect 1595 119 1599 123
rect 1601 119 1605 123
rect 1607 119 1611 123
rect 1613 119 1617 123
rect 1577 107 1581 111
rect 1583 107 1587 111
rect 1589 107 1593 111
rect 1595 107 1599 111
rect 1601 107 1605 111
rect 1607 107 1611 111
rect 1613 107 1617 111
rect 1443 92 1447 101
rect 1449 92 1453 101
rect 1455 92 1459 101
rect 1461 92 1465 101
rect 1467 92 1471 101
rect 1473 92 1477 101
rect 1479 92 1483 101
rect 1443 86 1447 90
rect 1449 86 1453 90
rect 1455 86 1459 90
rect 1461 86 1465 90
rect 1467 86 1471 90
rect 1473 86 1477 90
rect 1479 86 1483 90
rect 1443 80 1447 84
rect 1449 80 1453 84
rect 1455 80 1459 84
rect 1461 80 1465 84
rect 1467 80 1471 84
rect 1473 80 1477 84
rect 1479 80 1483 84
rect 1443 74 1447 78
rect 1449 74 1453 78
rect 1455 74 1459 78
rect 1461 74 1465 78
rect 1467 74 1471 78
rect 1473 74 1477 78
rect 1479 74 1483 78
rect 1443 63 1447 72
rect 1449 63 1453 72
rect 1455 63 1459 72
rect 1461 63 1465 72
rect 1467 63 1471 72
rect 1473 63 1477 72
rect 1479 63 1483 72
rect 1443 0 1447 4
rect 1449 0 1453 4
rect 1455 0 1459 4
rect 1461 0 1465 4
rect 1467 0 1471 4
rect 1473 0 1477 4
rect 1479 0 1483 4
rect 1526 53 1530 57
rect 1536 53 1540 57
rect 1487 44 1491 48
rect 1493 44 1497 48
rect 1499 44 1503 48
rect 1505 44 1509 48
rect 1511 44 1515 48
rect 1517 44 1521 48
rect 1523 44 1527 48
rect 1487 32 1491 36
rect 1493 32 1497 36
rect 1499 32 1503 36
rect 1505 32 1509 36
rect 1511 32 1515 36
rect 1517 32 1521 36
rect 1523 32 1527 36
rect 1487 26 1491 30
rect 1493 26 1497 30
rect 1499 26 1503 30
rect 1505 26 1509 30
rect 1511 26 1515 30
rect 1517 26 1521 30
rect 1523 26 1527 30
rect 1493 14 1497 18
rect 1499 14 1503 18
rect 1505 14 1509 18
rect 1511 14 1515 18
rect 1517 14 1521 18
rect 1523 14 1527 18
rect 1487 0 1491 4
rect 1493 0 1497 4
rect 1499 0 1503 4
rect 1505 0 1509 4
rect 1511 0 1515 4
rect 1517 0 1521 4
rect 1523 0 1527 4
rect 1531 0 1540 4
rect 1564 53 1568 57
rect 1574 53 1578 57
rect 1564 0 1573 4
rect 1577 44 1581 48
rect 1583 44 1587 48
rect 1589 44 1593 48
rect 1595 44 1599 48
rect 1601 44 1605 48
rect 1607 44 1611 48
rect 1613 44 1617 48
rect 1577 32 1581 36
rect 1583 32 1587 36
rect 1589 32 1593 36
rect 1595 32 1599 36
rect 1601 32 1605 36
rect 1607 32 1611 36
rect 1613 32 1617 36
rect 1577 26 1581 30
rect 1583 26 1587 30
rect 1589 26 1593 30
rect 1595 26 1599 30
rect 1601 26 1605 30
rect 1607 26 1611 30
rect 1613 26 1617 30
rect 1577 14 1581 18
rect 1583 14 1587 18
rect 1589 14 1593 18
rect 1595 14 1599 18
rect 1601 14 1605 18
rect 1607 14 1611 18
rect 1577 0 1581 4
rect 1583 0 1587 4
rect 1589 0 1593 4
rect 1595 0 1599 4
rect 1601 0 1605 4
rect 1607 0 1611 4
rect 1613 0 1617 4
rect 1621 92 1625 101
rect 1627 92 1631 101
rect 1633 92 1637 101
rect 1639 92 1643 101
rect 1645 92 1649 101
rect 1651 92 1655 101
rect 1657 92 1661 101
rect 1621 86 1625 90
rect 1627 86 1631 90
rect 1633 86 1637 90
rect 1639 86 1643 90
rect 1645 86 1649 90
rect 1651 86 1655 90
rect 1657 86 1661 90
rect 1621 80 1625 84
rect 1627 80 1631 84
rect 1633 80 1637 84
rect 1639 80 1643 84
rect 1645 80 1649 84
rect 1651 80 1655 84
rect 1657 80 1661 84
rect 1621 74 1625 78
rect 1627 74 1631 78
rect 1633 74 1637 78
rect 1639 74 1643 78
rect 1645 74 1649 78
rect 1651 74 1655 78
rect 1657 74 1661 78
rect 1621 63 1625 72
rect 1627 63 1631 72
rect 1633 63 1637 72
rect 1639 63 1643 72
rect 1645 63 1649 72
rect 1651 63 1655 72
rect 1657 63 1661 72
rect 1621 0 1625 4
rect 1627 0 1631 4
rect 1633 0 1637 4
rect 1639 0 1643 4
rect 1645 0 1649 4
rect 1651 0 1655 4
rect 1657 0 1661 4
rect 1967 131 1971 135
rect 1973 131 1977 135
rect 1979 131 1983 135
rect 1985 131 1989 135
rect 1991 131 1995 135
rect 1997 131 2001 135
rect 1961 119 1965 123
rect 1967 119 1971 123
rect 1973 119 1977 123
rect 1979 119 1983 123
rect 1985 119 1989 123
rect 1991 119 1995 123
rect 1997 119 2001 123
rect 1961 107 1965 111
rect 1967 107 1971 111
rect 1973 107 1977 111
rect 1979 107 1983 111
rect 1985 107 1989 111
rect 1991 107 1995 111
rect 1997 107 2001 111
rect 2051 131 2055 135
rect 2057 131 2061 135
rect 2063 131 2067 135
rect 2069 131 2073 135
rect 2075 131 2079 135
rect 2081 131 2085 135
rect 2051 119 2055 123
rect 2057 119 2061 123
rect 2063 119 2067 123
rect 2069 119 2073 123
rect 2075 119 2079 123
rect 2081 119 2085 123
rect 2087 119 2091 123
rect 2051 107 2055 111
rect 2057 107 2061 111
rect 2063 107 2067 111
rect 2069 107 2073 111
rect 2075 107 2079 111
rect 2081 107 2085 111
rect 2087 107 2091 111
rect 1917 92 1921 101
rect 1923 92 1927 101
rect 1929 92 1933 101
rect 1935 92 1939 101
rect 1941 92 1945 101
rect 1947 92 1951 101
rect 1953 92 1957 101
rect 1917 86 1921 90
rect 1923 86 1927 90
rect 1929 86 1933 90
rect 1935 86 1939 90
rect 1941 86 1945 90
rect 1947 86 1951 90
rect 1953 86 1957 90
rect 1917 80 1921 84
rect 1923 80 1927 84
rect 1929 80 1933 84
rect 1935 80 1939 84
rect 1941 80 1945 84
rect 1947 80 1951 84
rect 1953 80 1957 84
rect 1917 74 1921 78
rect 1923 74 1927 78
rect 1929 74 1933 78
rect 1935 74 1939 78
rect 1941 74 1945 78
rect 1947 74 1951 78
rect 1953 74 1957 78
rect 1917 63 1921 72
rect 1923 63 1927 72
rect 1929 63 1933 72
rect 1935 63 1939 72
rect 1941 63 1945 72
rect 1947 63 1951 72
rect 1953 63 1957 72
rect 1917 0 1921 4
rect 1923 0 1927 4
rect 1929 0 1933 4
rect 1935 0 1939 4
rect 1941 0 1945 4
rect 1947 0 1951 4
rect 1953 0 1957 4
rect 2000 53 2004 57
rect 2010 53 2014 57
rect 1961 44 1965 48
rect 1967 44 1971 48
rect 1973 44 1977 48
rect 1979 44 1983 48
rect 1985 44 1989 48
rect 1991 44 1995 48
rect 1997 44 2001 48
rect 1961 32 1965 36
rect 1967 32 1971 36
rect 1973 32 1977 36
rect 1979 32 1983 36
rect 1985 32 1989 36
rect 1991 32 1995 36
rect 1997 32 2001 36
rect 1961 26 1965 30
rect 1967 26 1971 30
rect 1973 26 1977 30
rect 1979 26 1983 30
rect 1985 26 1989 30
rect 1991 26 1995 30
rect 1997 26 2001 30
rect 1967 14 1971 18
rect 1973 14 1977 18
rect 1979 14 1983 18
rect 1985 14 1989 18
rect 1991 14 1995 18
rect 1997 14 2001 18
rect 1961 0 1965 4
rect 1967 0 1971 4
rect 1973 0 1977 4
rect 1979 0 1983 4
rect 1985 0 1989 4
rect 1991 0 1995 4
rect 1997 0 2001 4
rect 2005 0 2014 4
rect 2038 53 2042 57
rect 2048 53 2052 57
rect 2038 0 2047 4
rect 2051 44 2055 48
rect 2057 44 2061 48
rect 2063 44 2067 48
rect 2069 44 2073 48
rect 2075 44 2079 48
rect 2081 44 2085 48
rect 2087 44 2091 48
rect 2051 32 2055 36
rect 2057 32 2061 36
rect 2063 32 2067 36
rect 2069 32 2073 36
rect 2075 32 2079 36
rect 2081 32 2085 36
rect 2087 32 2091 36
rect 2051 26 2055 30
rect 2057 26 2061 30
rect 2063 26 2067 30
rect 2069 26 2073 30
rect 2075 26 2079 30
rect 2081 26 2085 30
rect 2087 26 2091 30
rect 2051 14 2055 18
rect 2057 14 2061 18
rect 2063 14 2067 18
rect 2069 14 2073 18
rect 2075 14 2079 18
rect 2081 14 2085 18
rect 2051 0 2055 4
rect 2057 0 2061 4
rect 2063 0 2067 4
rect 2069 0 2073 4
rect 2075 0 2079 4
rect 2081 0 2085 4
rect 2087 0 2091 4
rect 2095 92 2099 101
rect 2101 92 2105 101
rect 2107 92 2111 101
rect 2113 92 2117 101
rect 2119 92 2123 101
rect 2125 92 2129 101
rect 2131 92 2135 101
rect 2095 86 2099 90
rect 2101 86 2105 90
rect 2107 86 2111 90
rect 2113 86 2117 90
rect 2119 86 2123 90
rect 2125 86 2129 90
rect 2131 86 2135 90
rect 2095 80 2099 84
rect 2101 80 2105 84
rect 2107 80 2111 84
rect 2113 80 2117 84
rect 2119 80 2123 84
rect 2125 80 2129 84
rect 2131 80 2135 84
rect 2095 74 2099 78
rect 2101 74 2105 78
rect 2107 74 2111 78
rect 2113 74 2117 78
rect 2119 74 2123 78
rect 2125 74 2129 78
rect 2131 74 2135 78
rect 2095 63 2099 72
rect 2101 63 2105 72
rect 2107 63 2111 72
rect 2113 63 2117 72
rect 2119 63 2123 72
rect 2125 63 2129 72
rect 2131 63 2135 72
rect 2095 0 2099 4
rect 2101 0 2105 4
rect 2107 0 2111 4
rect 2113 0 2117 4
rect 2119 0 2123 4
rect 2125 0 2129 4
rect 2131 0 2135 4
rect 2441 131 2445 135
rect 2447 131 2451 135
rect 2453 131 2457 135
rect 2459 131 2463 135
rect 2465 131 2469 135
rect 2471 131 2475 135
rect 2435 119 2439 123
rect 2441 119 2445 123
rect 2447 119 2451 123
rect 2453 119 2457 123
rect 2459 119 2463 123
rect 2465 119 2469 123
rect 2471 119 2475 123
rect 2435 107 2439 111
rect 2441 107 2445 111
rect 2447 107 2451 111
rect 2453 107 2457 111
rect 2459 107 2463 111
rect 2465 107 2469 111
rect 2471 107 2475 111
rect 2525 131 2529 135
rect 2531 131 2535 135
rect 2537 131 2541 135
rect 2543 131 2547 135
rect 2549 131 2553 135
rect 2555 131 2559 135
rect 2525 119 2529 123
rect 2531 119 2535 123
rect 2537 119 2541 123
rect 2543 119 2547 123
rect 2549 119 2553 123
rect 2555 119 2559 123
rect 2561 119 2565 123
rect 2525 107 2529 111
rect 2531 107 2535 111
rect 2537 107 2541 111
rect 2543 107 2547 111
rect 2549 107 2553 111
rect 2555 107 2559 111
rect 2561 107 2565 111
rect 2391 92 2395 101
rect 2397 92 2401 101
rect 2403 92 2407 101
rect 2409 92 2413 101
rect 2415 92 2419 101
rect 2421 92 2425 101
rect 2427 92 2431 101
rect 2391 86 2395 90
rect 2397 86 2401 90
rect 2403 86 2407 90
rect 2409 86 2413 90
rect 2415 86 2419 90
rect 2421 86 2425 90
rect 2427 86 2431 90
rect 2391 80 2395 84
rect 2397 80 2401 84
rect 2403 80 2407 84
rect 2409 80 2413 84
rect 2415 80 2419 84
rect 2421 80 2425 84
rect 2427 80 2431 84
rect 2391 74 2395 78
rect 2397 74 2401 78
rect 2403 74 2407 78
rect 2409 74 2413 78
rect 2415 74 2419 78
rect 2421 74 2425 78
rect 2427 74 2431 78
rect 2391 63 2395 72
rect 2397 63 2401 72
rect 2403 63 2407 72
rect 2409 63 2413 72
rect 2415 63 2419 72
rect 2421 63 2425 72
rect 2427 63 2431 72
rect 2391 0 2395 4
rect 2397 0 2401 4
rect 2403 0 2407 4
rect 2409 0 2413 4
rect 2415 0 2419 4
rect 2421 0 2425 4
rect 2427 0 2431 4
rect 2474 53 2478 57
rect 2484 53 2488 57
rect 2435 44 2439 48
rect 2441 44 2445 48
rect 2447 44 2451 48
rect 2453 44 2457 48
rect 2459 44 2463 48
rect 2465 44 2469 48
rect 2471 44 2475 48
rect 2435 32 2439 36
rect 2441 32 2445 36
rect 2447 32 2451 36
rect 2453 32 2457 36
rect 2459 32 2463 36
rect 2465 32 2469 36
rect 2471 32 2475 36
rect 2435 26 2439 30
rect 2441 26 2445 30
rect 2447 26 2451 30
rect 2453 26 2457 30
rect 2459 26 2463 30
rect 2465 26 2469 30
rect 2471 26 2475 30
rect 2441 14 2445 18
rect 2447 14 2451 18
rect 2453 14 2457 18
rect 2459 14 2463 18
rect 2465 14 2469 18
rect 2471 14 2475 18
rect 2435 0 2439 4
rect 2441 0 2445 4
rect 2447 0 2451 4
rect 2453 0 2457 4
rect 2459 0 2463 4
rect 2465 0 2469 4
rect 2471 0 2475 4
rect 2479 0 2488 4
rect 2512 53 2516 57
rect 2522 53 2526 57
rect 2512 0 2521 4
rect 2525 44 2529 48
rect 2531 44 2535 48
rect 2537 44 2541 48
rect 2543 44 2547 48
rect 2549 44 2553 48
rect 2555 44 2559 48
rect 2561 44 2565 48
rect 2525 32 2529 36
rect 2531 32 2535 36
rect 2537 32 2541 36
rect 2543 32 2547 36
rect 2549 32 2553 36
rect 2555 32 2559 36
rect 2561 32 2565 36
rect 2525 26 2529 30
rect 2531 26 2535 30
rect 2537 26 2541 30
rect 2543 26 2547 30
rect 2549 26 2553 30
rect 2555 26 2559 30
rect 2561 26 2565 30
rect 2525 14 2529 18
rect 2531 14 2535 18
rect 2537 14 2541 18
rect 2543 14 2547 18
rect 2549 14 2553 18
rect 2555 14 2559 18
rect 2525 0 2529 4
rect 2531 0 2535 4
rect 2537 0 2541 4
rect 2543 0 2547 4
rect 2549 0 2553 4
rect 2555 0 2559 4
rect 2561 0 2565 4
rect 2569 92 2573 101
rect 2575 92 2579 101
rect 2581 92 2585 101
rect 2587 92 2591 101
rect 2593 92 2597 101
rect 2599 92 2603 101
rect 2605 92 2609 101
rect 2569 86 2573 90
rect 2575 86 2579 90
rect 2581 86 2585 90
rect 2587 86 2591 90
rect 2593 86 2597 90
rect 2599 86 2603 90
rect 2605 86 2609 90
rect 2569 80 2573 84
rect 2575 80 2579 84
rect 2581 80 2585 84
rect 2587 80 2591 84
rect 2593 80 2597 84
rect 2599 80 2603 84
rect 2605 80 2609 84
rect 2569 74 2573 78
rect 2575 74 2579 78
rect 2581 74 2585 78
rect 2587 74 2591 78
rect 2593 74 2597 78
rect 2599 74 2603 78
rect 2605 74 2609 78
rect 2569 63 2573 72
rect 2575 63 2579 72
rect 2581 63 2585 72
rect 2587 63 2591 72
rect 2593 63 2597 72
rect 2599 63 2603 72
rect 2605 63 2609 72
rect 2569 0 2573 4
rect 2575 0 2579 4
rect 2581 0 2585 4
rect 2587 0 2591 4
rect 2593 0 2597 4
rect 2599 0 2603 4
rect 2605 0 2609 4
rect 2915 131 2919 135
rect 2921 131 2925 135
rect 2927 131 2931 135
rect 2933 131 2937 135
rect 2939 131 2943 135
rect 2945 131 2949 135
rect 2909 119 2913 123
rect 2915 119 2919 123
rect 2921 119 2925 123
rect 2927 119 2931 123
rect 2933 119 2937 123
rect 2939 119 2943 123
rect 2945 119 2949 123
rect 2909 107 2913 111
rect 2915 107 2919 111
rect 2921 107 2925 111
rect 2927 107 2931 111
rect 2933 107 2937 111
rect 2939 107 2943 111
rect 2945 107 2949 111
rect 2999 131 3003 135
rect 3005 131 3009 135
rect 3011 131 3015 135
rect 3017 131 3021 135
rect 3023 131 3027 135
rect 3029 131 3033 135
rect 2999 119 3003 123
rect 3005 119 3009 123
rect 3011 119 3015 123
rect 3017 119 3021 123
rect 3023 119 3027 123
rect 3029 119 3033 123
rect 3035 119 3039 123
rect 2999 107 3003 111
rect 3005 107 3009 111
rect 3011 107 3015 111
rect 3017 107 3021 111
rect 3023 107 3027 111
rect 3029 107 3033 111
rect 3035 107 3039 111
rect 2865 92 2869 101
rect 2871 92 2875 101
rect 2877 92 2881 101
rect 2883 92 2887 101
rect 2889 92 2893 101
rect 2895 92 2899 101
rect 2901 92 2905 101
rect 2865 86 2869 90
rect 2871 86 2875 90
rect 2877 86 2881 90
rect 2883 86 2887 90
rect 2889 86 2893 90
rect 2895 86 2899 90
rect 2901 86 2905 90
rect 2865 80 2869 84
rect 2871 80 2875 84
rect 2877 80 2881 84
rect 2883 80 2887 84
rect 2889 80 2893 84
rect 2895 80 2899 84
rect 2901 80 2905 84
rect 2865 74 2869 78
rect 2871 74 2875 78
rect 2877 74 2881 78
rect 2883 74 2887 78
rect 2889 74 2893 78
rect 2895 74 2899 78
rect 2901 74 2905 78
rect 2865 63 2869 72
rect 2871 63 2875 72
rect 2877 63 2881 72
rect 2883 63 2887 72
rect 2889 63 2893 72
rect 2895 63 2899 72
rect 2901 63 2905 72
rect 2865 0 2869 4
rect 2871 0 2875 4
rect 2877 0 2881 4
rect 2883 0 2887 4
rect 2889 0 2893 4
rect 2895 0 2899 4
rect 2901 0 2905 4
rect 2948 53 2952 57
rect 2958 53 2962 57
rect 2909 44 2913 48
rect 2915 44 2919 48
rect 2921 44 2925 48
rect 2927 44 2931 48
rect 2933 44 2937 48
rect 2939 44 2943 48
rect 2945 44 2949 48
rect 2909 32 2913 36
rect 2915 32 2919 36
rect 2921 32 2925 36
rect 2927 32 2931 36
rect 2933 32 2937 36
rect 2939 32 2943 36
rect 2945 32 2949 36
rect 2909 26 2913 30
rect 2915 26 2919 30
rect 2921 26 2925 30
rect 2927 26 2931 30
rect 2933 26 2937 30
rect 2939 26 2943 30
rect 2945 26 2949 30
rect 2915 14 2919 18
rect 2921 14 2925 18
rect 2927 14 2931 18
rect 2933 14 2937 18
rect 2939 14 2943 18
rect 2945 14 2949 18
rect 2909 0 2913 4
rect 2915 0 2919 4
rect 2921 0 2925 4
rect 2927 0 2931 4
rect 2933 0 2937 4
rect 2939 0 2943 4
rect 2945 0 2949 4
rect 2953 0 2962 4
rect 2986 53 2990 57
rect 2996 53 3000 57
rect 2986 0 2995 4
rect 2999 44 3003 48
rect 3005 44 3009 48
rect 3011 44 3015 48
rect 3017 44 3021 48
rect 3023 44 3027 48
rect 3029 44 3033 48
rect 3035 44 3039 48
rect 2999 32 3003 36
rect 3005 32 3009 36
rect 3011 32 3015 36
rect 3017 32 3021 36
rect 3023 32 3027 36
rect 3029 32 3033 36
rect 3035 32 3039 36
rect 2999 26 3003 30
rect 3005 26 3009 30
rect 3011 26 3015 30
rect 3017 26 3021 30
rect 3023 26 3027 30
rect 3029 26 3033 30
rect 3035 26 3039 30
rect 2999 14 3003 18
rect 3005 14 3009 18
rect 3011 14 3015 18
rect 3017 14 3021 18
rect 3023 14 3027 18
rect 3029 14 3033 18
rect 2999 0 3003 4
rect 3005 0 3009 4
rect 3011 0 3015 4
rect 3017 0 3021 4
rect 3023 0 3027 4
rect 3029 0 3033 4
rect 3035 0 3039 4
rect 3043 92 3047 101
rect 3049 92 3053 101
rect 3055 92 3059 101
rect 3061 92 3065 101
rect 3067 92 3071 101
rect 3073 92 3077 101
rect 3079 92 3083 101
rect 3043 86 3047 90
rect 3049 86 3053 90
rect 3055 86 3059 90
rect 3061 86 3065 90
rect 3067 86 3071 90
rect 3073 86 3077 90
rect 3079 86 3083 90
rect 3043 80 3047 84
rect 3049 80 3053 84
rect 3055 80 3059 84
rect 3061 80 3065 84
rect 3067 80 3071 84
rect 3073 80 3077 84
rect 3079 80 3083 84
rect 3043 74 3047 78
rect 3049 74 3053 78
rect 3055 74 3059 78
rect 3061 74 3065 78
rect 3067 74 3071 78
rect 3073 74 3077 78
rect 3079 74 3083 78
rect 3043 63 3047 72
rect 3049 63 3053 72
rect 3055 63 3059 72
rect 3061 63 3065 72
rect 3067 63 3071 72
rect 3073 63 3077 72
rect 3079 63 3083 72
rect 3043 0 3047 4
rect 3049 0 3053 4
rect 3055 0 3059 4
rect 3061 0 3065 4
rect 3067 0 3071 4
rect 3073 0 3077 4
rect 3079 0 3083 4
rect 3389 131 3393 135
rect 3395 131 3399 135
rect 3401 131 3405 135
rect 3407 131 3411 135
rect 3413 131 3417 135
rect 3419 131 3423 135
rect 3383 119 3387 123
rect 3389 119 3393 123
rect 3395 119 3399 123
rect 3401 119 3405 123
rect 3407 119 3411 123
rect 3413 119 3417 123
rect 3419 119 3423 123
rect 3383 107 3387 111
rect 3389 107 3393 111
rect 3395 107 3399 111
rect 3401 107 3405 111
rect 3407 107 3411 111
rect 3413 107 3417 111
rect 3419 107 3423 111
rect 3473 131 3477 135
rect 3479 131 3483 135
rect 3485 131 3489 135
rect 3491 131 3495 135
rect 3497 131 3501 135
rect 3503 131 3507 135
rect 3473 119 3477 123
rect 3479 119 3483 123
rect 3485 119 3489 123
rect 3491 119 3495 123
rect 3497 119 3501 123
rect 3503 119 3507 123
rect 3509 119 3513 123
rect 3473 107 3477 111
rect 3479 107 3483 111
rect 3485 107 3489 111
rect 3491 107 3495 111
rect 3497 107 3501 111
rect 3503 107 3507 111
rect 3509 107 3513 111
rect 3339 92 3343 101
rect 3345 92 3349 101
rect 3351 92 3355 101
rect 3357 92 3361 101
rect 3363 92 3367 101
rect 3369 92 3373 101
rect 3375 92 3379 101
rect 3339 86 3343 90
rect 3345 86 3349 90
rect 3351 86 3355 90
rect 3357 86 3361 90
rect 3363 86 3367 90
rect 3369 86 3373 90
rect 3375 86 3379 90
rect 3339 80 3343 84
rect 3345 80 3349 84
rect 3351 80 3355 84
rect 3357 80 3361 84
rect 3363 80 3367 84
rect 3369 80 3373 84
rect 3375 80 3379 84
rect 3339 74 3343 78
rect 3345 74 3349 78
rect 3351 74 3355 78
rect 3357 74 3361 78
rect 3363 74 3367 78
rect 3369 74 3373 78
rect 3375 74 3379 78
rect 3339 63 3343 72
rect 3345 63 3349 72
rect 3351 63 3355 72
rect 3357 63 3361 72
rect 3363 63 3367 72
rect 3369 63 3373 72
rect 3375 63 3379 72
rect 3339 0 3343 4
rect 3345 0 3349 4
rect 3351 0 3355 4
rect 3357 0 3361 4
rect 3363 0 3367 4
rect 3369 0 3373 4
rect 3375 0 3379 4
rect 3422 53 3426 57
rect 3432 53 3436 57
rect 3383 44 3387 48
rect 3389 44 3393 48
rect 3395 44 3399 48
rect 3401 44 3405 48
rect 3407 44 3411 48
rect 3413 44 3417 48
rect 3419 44 3423 48
rect 3383 32 3387 36
rect 3389 32 3393 36
rect 3395 32 3399 36
rect 3401 32 3405 36
rect 3407 32 3411 36
rect 3413 32 3417 36
rect 3419 32 3423 36
rect 3383 26 3387 30
rect 3389 26 3393 30
rect 3395 26 3399 30
rect 3401 26 3405 30
rect 3407 26 3411 30
rect 3413 26 3417 30
rect 3419 26 3423 30
rect 3389 14 3393 18
rect 3395 14 3399 18
rect 3401 14 3405 18
rect 3407 14 3411 18
rect 3413 14 3417 18
rect 3419 14 3423 18
rect 3383 0 3387 4
rect 3389 0 3393 4
rect 3395 0 3399 4
rect 3401 0 3405 4
rect 3407 0 3411 4
rect 3413 0 3417 4
rect 3419 0 3423 4
rect 3427 0 3436 4
rect 3460 53 3464 57
rect 3470 53 3474 57
rect 3460 0 3469 4
rect 3473 44 3477 48
rect 3479 44 3483 48
rect 3485 44 3489 48
rect 3491 44 3495 48
rect 3497 44 3501 48
rect 3503 44 3507 48
rect 3509 44 3513 48
rect 3473 32 3477 36
rect 3479 32 3483 36
rect 3485 32 3489 36
rect 3491 32 3495 36
rect 3497 32 3501 36
rect 3503 32 3507 36
rect 3509 32 3513 36
rect 3473 26 3477 30
rect 3479 26 3483 30
rect 3485 26 3489 30
rect 3491 26 3495 30
rect 3497 26 3501 30
rect 3503 26 3507 30
rect 3509 26 3513 30
rect 3473 14 3477 18
rect 3479 14 3483 18
rect 3485 14 3489 18
rect 3491 14 3495 18
rect 3497 14 3501 18
rect 3503 14 3507 18
rect 3473 0 3477 4
rect 3479 0 3483 4
rect 3485 0 3489 4
rect 3491 0 3495 4
rect 3497 0 3501 4
rect 3503 0 3507 4
rect 3509 0 3513 4
rect 3517 92 3521 101
rect 3523 92 3527 101
rect 3529 92 3533 101
rect 3535 92 3539 101
rect 3541 92 3545 101
rect 3547 92 3551 101
rect 3553 92 3557 101
rect 3517 86 3521 90
rect 3523 86 3527 90
rect 3529 86 3533 90
rect 3535 86 3539 90
rect 3541 86 3545 90
rect 3547 86 3551 90
rect 3553 86 3557 90
rect 3517 80 3521 84
rect 3523 80 3527 84
rect 3529 80 3533 84
rect 3535 80 3539 84
rect 3541 80 3545 84
rect 3547 80 3551 84
rect 3553 80 3557 84
rect 3517 74 3521 78
rect 3523 74 3527 78
rect 3529 74 3533 78
rect 3535 74 3539 78
rect 3541 74 3545 78
rect 3547 74 3551 78
rect 3553 74 3557 78
rect 3517 63 3521 72
rect 3523 63 3527 72
rect 3529 63 3533 72
rect 3535 63 3539 72
rect 3541 63 3545 72
rect 3547 63 3551 72
rect 3553 63 3557 72
rect 3517 0 3521 4
rect 3523 0 3527 4
rect 3529 0 3533 4
rect 3535 0 3539 4
rect 3541 0 3545 4
rect 3547 0 3551 4
rect 3553 0 3557 4
rect 3863 131 3867 135
rect 3869 131 3873 135
rect 3875 131 3879 135
rect 3881 131 3885 135
rect 3887 131 3891 135
rect 3893 131 3897 135
rect 3857 119 3861 123
rect 3863 119 3867 123
rect 3869 119 3873 123
rect 3875 119 3879 123
rect 3881 119 3885 123
rect 3887 119 3891 123
rect 3893 119 3897 123
rect 3857 107 3861 111
rect 3863 107 3867 111
rect 3869 107 3873 111
rect 3875 107 3879 111
rect 3881 107 3885 111
rect 3887 107 3891 111
rect 3893 107 3897 111
rect 3947 131 3951 135
rect 3953 131 3957 135
rect 3959 131 3963 135
rect 3965 131 3969 135
rect 3971 131 3975 135
rect 3977 131 3981 135
rect 3947 119 3951 123
rect 3953 119 3957 123
rect 3959 119 3963 123
rect 3965 119 3969 123
rect 3971 119 3975 123
rect 3977 119 3981 123
rect 3983 119 3987 123
rect 3947 107 3951 111
rect 3953 107 3957 111
rect 3959 107 3963 111
rect 3965 107 3969 111
rect 3971 107 3975 111
rect 3977 107 3981 111
rect 3983 107 3987 111
rect 3813 92 3817 101
rect 3819 92 3823 101
rect 3825 92 3829 101
rect 3831 92 3835 101
rect 3837 92 3841 101
rect 3843 92 3847 101
rect 3849 92 3853 101
rect 3813 86 3817 90
rect 3819 86 3823 90
rect 3825 86 3829 90
rect 3831 86 3835 90
rect 3837 86 3841 90
rect 3843 86 3847 90
rect 3849 86 3853 90
rect 3813 80 3817 84
rect 3819 80 3823 84
rect 3825 80 3829 84
rect 3831 80 3835 84
rect 3837 80 3841 84
rect 3843 80 3847 84
rect 3849 80 3853 84
rect 3813 74 3817 78
rect 3819 74 3823 78
rect 3825 74 3829 78
rect 3831 74 3835 78
rect 3837 74 3841 78
rect 3843 74 3847 78
rect 3849 74 3853 78
rect 3813 63 3817 72
rect 3819 63 3823 72
rect 3825 63 3829 72
rect 3831 63 3835 72
rect 3837 63 3841 72
rect 3843 63 3847 72
rect 3849 63 3853 72
rect 3813 0 3817 4
rect 3819 0 3823 4
rect 3825 0 3829 4
rect 3831 0 3835 4
rect 3837 0 3841 4
rect 3843 0 3847 4
rect 3849 0 3853 4
rect 3896 53 3900 57
rect 3906 53 3910 57
rect 3857 44 3861 48
rect 3863 44 3867 48
rect 3869 44 3873 48
rect 3875 44 3879 48
rect 3881 44 3885 48
rect 3887 44 3891 48
rect 3893 44 3897 48
rect 3857 32 3861 36
rect 3863 32 3867 36
rect 3869 32 3873 36
rect 3875 32 3879 36
rect 3881 32 3885 36
rect 3887 32 3891 36
rect 3893 32 3897 36
rect 3857 26 3861 30
rect 3863 26 3867 30
rect 3869 26 3873 30
rect 3875 26 3879 30
rect 3881 26 3885 30
rect 3887 26 3891 30
rect 3893 26 3897 30
rect 3863 14 3867 18
rect 3869 14 3873 18
rect 3875 14 3879 18
rect 3881 14 3885 18
rect 3887 14 3891 18
rect 3893 14 3897 18
rect 3857 0 3861 4
rect 3863 0 3867 4
rect 3869 0 3873 4
rect 3875 0 3879 4
rect 3881 0 3885 4
rect 3887 0 3891 4
rect 3893 0 3897 4
rect 3901 0 3910 4
rect 3934 53 3938 57
rect 3944 53 3948 57
rect 3934 0 3943 4
rect 3947 44 3951 48
rect 3953 44 3957 48
rect 3959 44 3963 48
rect 3965 44 3969 48
rect 3971 44 3975 48
rect 3977 44 3981 48
rect 3983 44 3987 48
rect 3947 32 3951 36
rect 3953 32 3957 36
rect 3959 32 3963 36
rect 3965 32 3969 36
rect 3971 32 3975 36
rect 3977 32 3981 36
rect 3983 32 3987 36
rect 3947 26 3951 30
rect 3953 26 3957 30
rect 3959 26 3963 30
rect 3965 26 3969 30
rect 3971 26 3975 30
rect 3977 26 3981 30
rect 3983 26 3987 30
rect 3947 14 3951 18
rect 3953 14 3957 18
rect 3959 14 3963 18
rect 3965 14 3969 18
rect 3971 14 3975 18
rect 3977 14 3981 18
rect 3947 0 3951 4
rect 3953 0 3957 4
rect 3959 0 3963 4
rect 3965 0 3969 4
rect 3971 0 3975 4
rect 3977 0 3981 4
rect 3983 0 3987 4
rect 3991 92 3995 101
rect 3997 92 4001 101
rect 4003 92 4007 101
rect 4009 92 4013 101
rect 4015 92 4019 101
rect 4021 92 4025 101
rect 4027 92 4031 101
rect 3991 86 3995 90
rect 3997 86 4001 90
rect 4003 86 4007 90
rect 4009 86 4013 90
rect 4015 86 4019 90
rect 4021 86 4025 90
rect 4027 86 4031 90
rect 3991 80 3995 84
rect 3997 80 4001 84
rect 4003 80 4007 84
rect 4009 80 4013 84
rect 4015 80 4019 84
rect 4021 80 4025 84
rect 4027 80 4031 84
rect 3991 74 3995 78
rect 3997 74 4001 78
rect 4003 74 4007 78
rect 4009 74 4013 78
rect 4015 74 4019 78
rect 4021 74 4025 78
rect 4027 74 4031 78
rect 3991 63 3995 72
rect 3997 63 4001 72
rect 4003 63 4007 72
rect 4009 63 4013 72
rect 4015 63 4019 72
rect 4021 63 4025 72
rect 4027 63 4031 72
rect 3991 0 3995 4
rect 3997 0 4001 4
rect 4003 0 4007 4
rect 4009 0 4013 4
rect 4015 0 4019 4
rect 4021 0 4025 4
rect 4027 0 4031 4
rect 4337 131 4341 135
rect 4343 131 4347 135
rect 4349 131 4353 135
rect 4355 131 4359 135
rect 4361 131 4365 135
rect 4367 131 4371 135
rect 4331 119 4335 123
rect 4337 119 4341 123
rect 4343 119 4347 123
rect 4349 119 4353 123
rect 4355 119 4359 123
rect 4361 119 4365 123
rect 4367 119 4371 123
rect 4331 107 4335 111
rect 4337 107 4341 111
rect 4343 107 4347 111
rect 4349 107 4353 111
rect 4355 107 4359 111
rect 4361 107 4365 111
rect 4367 107 4371 111
rect 4421 131 4425 135
rect 4427 131 4431 135
rect 4433 131 4437 135
rect 4439 131 4443 135
rect 4445 131 4449 135
rect 4451 131 4455 135
rect 4421 119 4425 123
rect 4427 119 4431 123
rect 4433 119 4437 123
rect 4439 119 4443 123
rect 4445 119 4449 123
rect 4451 119 4455 123
rect 4457 119 4461 123
rect 4421 107 4425 111
rect 4427 107 4431 111
rect 4433 107 4437 111
rect 4439 107 4443 111
rect 4445 107 4449 111
rect 4451 107 4455 111
rect 4457 107 4461 111
rect 4287 92 4291 101
rect 4293 92 4297 101
rect 4299 92 4303 101
rect 4305 92 4309 101
rect 4311 92 4315 101
rect 4317 92 4321 101
rect 4323 92 4327 101
rect 4287 86 4291 90
rect 4293 86 4297 90
rect 4299 86 4303 90
rect 4305 86 4309 90
rect 4311 86 4315 90
rect 4317 86 4321 90
rect 4323 86 4327 90
rect 4287 80 4291 84
rect 4293 80 4297 84
rect 4299 80 4303 84
rect 4305 80 4309 84
rect 4311 80 4315 84
rect 4317 80 4321 84
rect 4323 80 4327 84
rect 4287 74 4291 78
rect 4293 74 4297 78
rect 4299 74 4303 78
rect 4305 74 4309 78
rect 4311 74 4315 78
rect 4317 74 4321 78
rect 4323 74 4327 78
rect 4287 63 4291 72
rect 4293 63 4297 72
rect 4299 63 4303 72
rect 4305 63 4309 72
rect 4311 63 4315 72
rect 4317 63 4321 72
rect 4323 63 4327 72
rect 4287 0 4291 4
rect 4293 0 4297 4
rect 4299 0 4303 4
rect 4305 0 4309 4
rect 4311 0 4315 4
rect 4317 0 4321 4
rect 4323 0 4327 4
rect 4370 53 4374 57
rect 4380 53 4384 57
rect 4331 44 4335 48
rect 4337 44 4341 48
rect 4343 44 4347 48
rect 4349 44 4353 48
rect 4355 44 4359 48
rect 4361 44 4365 48
rect 4367 44 4371 48
rect 4331 32 4335 36
rect 4337 32 4341 36
rect 4343 32 4347 36
rect 4349 32 4353 36
rect 4355 32 4359 36
rect 4361 32 4365 36
rect 4367 32 4371 36
rect 4331 26 4335 30
rect 4337 26 4341 30
rect 4343 26 4347 30
rect 4349 26 4353 30
rect 4355 26 4359 30
rect 4361 26 4365 30
rect 4367 26 4371 30
rect 4337 14 4341 18
rect 4343 14 4347 18
rect 4349 14 4353 18
rect 4355 14 4359 18
rect 4361 14 4365 18
rect 4367 14 4371 18
rect 4331 0 4335 4
rect 4337 0 4341 4
rect 4343 0 4347 4
rect 4349 0 4353 4
rect 4355 0 4359 4
rect 4361 0 4365 4
rect 4367 0 4371 4
rect 4375 0 4384 4
rect 4408 53 4412 57
rect 4418 53 4422 57
rect 4465 92 4469 101
rect 4471 92 4475 101
rect 4477 92 4481 101
rect 4483 92 4487 101
rect 4489 92 4493 101
rect 4495 92 4499 101
rect 4501 92 4505 101
rect 4465 86 4469 90
rect 4471 86 4475 90
rect 4477 86 4481 90
rect 4483 86 4487 90
rect 4489 86 4493 90
rect 4495 86 4499 90
rect 4501 86 4505 90
rect 4465 80 4469 84
rect 4471 80 4475 84
rect 4477 80 4481 84
rect 4483 80 4487 84
rect 4489 80 4493 84
rect 4495 80 4499 84
rect 4501 80 4505 84
rect 4465 74 4469 78
rect 4471 74 4475 78
rect 4477 74 4481 78
rect 4483 74 4487 78
rect 4489 74 4493 78
rect 4495 74 4499 78
rect 4501 74 4505 78
rect 4465 63 4469 72
rect 4471 63 4475 72
rect 4477 63 4481 72
rect 4483 63 4487 72
rect 4489 63 4493 72
rect 4495 63 4499 72
rect 4501 63 4505 72
rect 4408 0 4417 4
rect 4421 44 4425 48
rect 4427 44 4431 48
rect 4433 44 4437 48
rect 4439 44 4443 48
rect 4445 44 4449 48
rect 4451 44 4455 48
rect 4457 44 4461 48
rect 4421 32 4425 36
rect 4427 32 4431 36
rect 4433 32 4437 36
rect 4439 32 4443 36
rect 4445 32 4449 36
rect 4451 32 4455 36
rect 4457 32 4461 36
rect 4421 26 4425 30
rect 4427 26 4431 30
rect 4433 26 4437 30
rect 4439 26 4443 30
rect 4445 26 4449 30
rect 4451 26 4455 30
rect 4457 26 4461 30
rect 4421 14 4425 18
rect 4427 14 4431 18
rect 4433 14 4437 18
rect 4439 14 4443 18
rect 4445 14 4449 18
rect 4451 14 4455 18
rect 4457 14 4461 18
rect 4421 0 4425 4
rect 4427 0 4431 4
rect 4433 0 4437 4
rect 4439 0 4443 4
rect 4445 0 4449 4
rect 4451 0 4455 4
rect 4457 0 4461 4
<< metal2 >>
rect 4643 499 4668 500
rect 4643 490 4644 499
rect 4653 490 4654 499
rect 4643 489 4668 490
rect 4642 180 4648 181
rect 4642 176 4643 180
rect 4647 176 4648 180
rect 4642 172 4648 176
rect 4642 168 4643 172
rect 4647 168 4648 172
rect 4642 164 4648 168
rect 4642 161 4643 164
rect 4618 160 4643 161
rect 4647 161 4648 164
rect 4674 180 4680 181
rect 4674 176 4675 180
rect 4679 176 4680 180
rect 4674 172 4680 176
rect 4674 168 4675 172
rect 4679 168 4680 172
rect 4674 164 4680 168
rect 4674 161 4675 164
rect 4647 160 4675 161
rect 4679 161 4680 164
rect 4698 180 4704 181
rect 4698 176 4699 180
rect 4703 176 4704 180
rect 4698 172 4704 176
rect 4698 168 4699 172
rect 4703 168 4704 172
rect 4698 164 4704 168
rect 4698 161 4699 164
rect 4679 160 4699 161
rect 4703 161 4704 164
rect 4730 180 4736 181
rect 4730 176 4731 180
rect 4735 176 4736 180
rect 4730 172 4736 176
rect 4730 168 4731 172
rect 4735 168 4736 172
rect 4730 164 4736 168
rect 4730 161 4731 164
rect 4703 160 4731 161
rect 4735 160 4736 164
rect 4618 156 4651 160
rect 4655 156 4659 160
rect 4663 156 4667 160
rect 4671 156 4707 160
rect 4711 156 4715 160
rect 4719 156 4723 160
rect 4727 156 4736 160
rect 4618 146 4736 156
rect 367 135 4633 146
rect 367 131 545 135
rect 549 131 551 135
rect 555 131 557 135
rect 561 131 563 135
rect 567 131 569 135
rect 573 131 575 135
rect 579 131 629 135
rect 633 131 635 135
rect 639 131 641 135
rect 645 131 647 135
rect 651 131 653 135
rect 657 131 659 135
rect 663 131 1019 135
rect 1023 131 1025 135
rect 1029 131 1031 135
rect 1035 131 1037 135
rect 1041 131 1043 135
rect 1047 131 1049 135
rect 1053 131 1103 135
rect 1107 131 1109 135
rect 1113 131 1115 135
rect 1119 131 1121 135
rect 1125 131 1127 135
rect 1131 131 1133 135
rect 1137 131 1493 135
rect 1497 131 1499 135
rect 1503 131 1505 135
rect 1509 131 1511 135
rect 1515 131 1517 135
rect 1521 131 1523 135
rect 1527 131 1577 135
rect 1581 131 1583 135
rect 1587 131 1589 135
rect 1593 131 1595 135
rect 1599 131 1601 135
rect 1605 131 1607 135
rect 1611 131 1967 135
rect 1971 131 1973 135
rect 1977 131 1979 135
rect 1983 131 1985 135
rect 1989 131 1991 135
rect 1995 131 1997 135
rect 2001 131 2051 135
rect 2055 131 2057 135
rect 2061 131 2063 135
rect 2067 131 2069 135
rect 2073 131 2075 135
rect 2079 131 2081 135
rect 2085 131 2441 135
rect 2445 131 2447 135
rect 2451 131 2453 135
rect 2457 131 2459 135
rect 2463 131 2465 135
rect 2469 131 2471 135
rect 2475 131 2525 135
rect 2529 131 2531 135
rect 2535 131 2537 135
rect 2541 131 2543 135
rect 2547 131 2549 135
rect 2553 131 2555 135
rect 2559 131 2915 135
rect 2919 131 2921 135
rect 2925 131 2927 135
rect 2931 131 2933 135
rect 2937 131 2939 135
rect 2943 131 2945 135
rect 2949 131 2999 135
rect 3003 131 3005 135
rect 3009 131 3011 135
rect 3015 131 3017 135
rect 3021 131 3023 135
rect 3027 131 3029 135
rect 3033 131 3389 135
rect 3393 131 3395 135
rect 3399 131 3401 135
rect 3405 131 3407 135
rect 3411 131 3413 135
rect 3417 131 3419 135
rect 3423 131 3473 135
rect 3477 131 3479 135
rect 3483 131 3485 135
rect 3489 131 3491 135
rect 3495 131 3497 135
rect 3501 131 3503 135
rect 3507 131 3863 135
rect 3867 131 3869 135
rect 3873 131 3875 135
rect 3879 131 3881 135
rect 3885 131 3887 135
rect 3891 131 3893 135
rect 3897 131 3947 135
rect 3951 131 3953 135
rect 3957 131 3959 135
rect 3963 131 3965 135
rect 3969 131 3971 135
rect 3975 131 3977 135
rect 3981 131 4337 135
rect 4341 131 4343 135
rect 4347 131 4349 135
rect 4353 131 4355 135
rect 4359 131 4361 135
rect 4365 131 4367 135
rect 4371 131 4421 135
rect 4425 131 4427 135
rect 4431 131 4433 135
rect 4437 131 4439 135
rect 4443 131 4445 135
rect 4449 131 4451 135
rect 4455 131 4633 135
rect 367 123 4633 131
rect 367 119 539 123
rect 543 119 545 123
rect 549 119 551 123
rect 555 119 557 123
rect 561 119 563 123
rect 567 119 569 123
rect 573 119 575 123
rect 579 119 629 123
rect 633 119 635 123
rect 639 119 641 123
rect 645 119 647 123
rect 651 119 653 123
rect 657 119 659 123
rect 663 119 665 123
rect 669 119 1013 123
rect 1017 119 1019 123
rect 1023 119 1025 123
rect 1029 119 1031 123
rect 1035 119 1037 123
rect 1041 119 1043 123
rect 1047 119 1049 123
rect 1053 119 1103 123
rect 1107 119 1109 123
rect 1113 119 1115 123
rect 1119 119 1121 123
rect 1125 119 1127 123
rect 1131 119 1133 123
rect 1137 119 1139 123
rect 1143 119 1487 123
rect 1491 119 1493 123
rect 1497 119 1499 123
rect 1503 119 1505 123
rect 1509 119 1511 123
rect 1515 119 1517 123
rect 1521 119 1523 123
rect 1527 119 1577 123
rect 1581 119 1583 123
rect 1587 119 1589 123
rect 1593 119 1595 123
rect 1599 119 1601 123
rect 1605 119 1607 123
rect 1611 119 1613 123
rect 1617 119 1961 123
rect 1965 119 1967 123
rect 1971 119 1973 123
rect 1977 119 1979 123
rect 1983 119 1985 123
rect 1989 119 1991 123
rect 1995 119 1997 123
rect 2001 119 2051 123
rect 2055 119 2057 123
rect 2061 119 2063 123
rect 2067 119 2069 123
rect 2073 119 2075 123
rect 2079 119 2081 123
rect 2085 119 2087 123
rect 2091 119 2435 123
rect 2439 119 2441 123
rect 2445 119 2447 123
rect 2451 119 2453 123
rect 2457 119 2459 123
rect 2463 119 2465 123
rect 2469 119 2471 123
rect 2475 119 2525 123
rect 2529 119 2531 123
rect 2535 119 2537 123
rect 2541 119 2543 123
rect 2547 119 2549 123
rect 2553 119 2555 123
rect 2559 119 2561 123
rect 2565 119 2909 123
rect 2913 119 2915 123
rect 2919 119 2921 123
rect 2925 119 2927 123
rect 2931 119 2933 123
rect 2937 119 2939 123
rect 2943 119 2945 123
rect 2949 119 2999 123
rect 3003 119 3005 123
rect 3009 119 3011 123
rect 3015 119 3017 123
rect 3021 119 3023 123
rect 3027 119 3029 123
rect 3033 119 3035 123
rect 3039 119 3383 123
rect 3387 119 3389 123
rect 3393 119 3395 123
rect 3399 119 3401 123
rect 3405 119 3407 123
rect 3411 119 3413 123
rect 3417 119 3419 123
rect 3423 119 3473 123
rect 3477 119 3479 123
rect 3483 119 3485 123
rect 3489 119 3491 123
rect 3495 119 3497 123
rect 3501 119 3503 123
rect 3507 119 3509 123
rect 3513 119 3857 123
rect 3861 119 3863 123
rect 3867 119 3869 123
rect 3873 119 3875 123
rect 3879 119 3881 123
rect 3885 119 3887 123
rect 3891 119 3893 123
rect 3897 119 3947 123
rect 3951 119 3953 123
rect 3957 119 3959 123
rect 3963 119 3965 123
rect 3969 119 3971 123
rect 3975 119 3977 123
rect 3981 119 3983 123
rect 3987 119 4331 123
rect 4335 119 4337 123
rect 4341 119 4343 123
rect 4347 119 4349 123
rect 4353 119 4355 123
rect 4359 119 4361 123
rect 4365 119 4367 123
rect 4371 119 4421 123
rect 4425 119 4427 123
rect 4431 119 4433 123
rect 4437 119 4439 123
rect 4443 119 4445 123
rect 4449 119 4451 123
rect 4455 119 4457 123
rect 4461 119 4633 123
rect 367 111 4633 119
rect 367 107 539 111
rect 543 107 545 111
rect 549 107 551 111
rect 555 107 557 111
rect 561 107 563 111
rect 567 107 569 111
rect 573 107 575 111
rect 579 107 629 111
rect 633 107 635 111
rect 639 107 641 111
rect 645 107 647 111
rect 651 107 653 111
rect 657 107 659 111
rect 663 107 665 111
rect 669 107 1013 111
rect 1017 107 1019 111
rect 1023 107 1025 111
rect 1029 107 1031 111
rect 1035 107 1037 111
rect 1041 107 1043 111
rect 1047 107 1049 111
rect 1053 107 1103 111
rect 1107 107 1109 111
rect 1113 107 1115 111
rect 1119 107 1121 111
rect 1125 107 1127 111
rect 1131 107 1133 111
rect 1137 107 1139 111
rect 1143 107 1487 111
rect 1491 107 1493 111
rect 1497 107 1499 111
rect 1503 107 1505 111
rect 1509 107 1511 111
rect 1515 107 1517 111
rect 1521 107 1523 111
rect 1527 107 1577 111
rect 1581 107 1583 111
rect 1587 107 1589 111
rect 1593 107 1595 111
rect 1599 107 1601 111
rect 1605 107 1607 111
rect 1611 107 1613 111
rect 1617 107 1961 111
rect 1965 107 1967 111
rect 1971 107 1973 111
rect 1977 107 1979 111
rect 1983 107 1985 111
rect 1989 107 1991 111
rect 1995 107 1997 111
rect 2001 107 2051 111
rect 2055 107 2057 111
rect 2061 107 2063 111
rect 2067 107 2069 111
rect 2073 107 2075 111
rect 2079 107 2081 111
rect 2085 107 2087 111
rect 2091 107 2435 111
rect 2439 107 2441 111
rect 2445 107 2447 111
rect 2451 107 2453 111
rect 2457 107 2459 111
rect 2463 107 2465 111
rect 2469 107 2471 111
rect 2475 107 2525 111
rect 2529 107 2531 111
rect 2535 107 2537 111
rect 2541 107 2543 111
rect 2547 107 2549 111
rect 2553 107 2555 111
rect 2559 107 2561 111
rect 2565 107 2909 111
rect 2913 107 2915 111
rect 2919 107 2921 111
rect 2925 107 2927 111
rect 2931 107 2933 111
rect 2937 107 2939 111
rect 2943 107 2945 111
rect 2949 107 2999 111
rect 3003 107 3005 111
rect 3009 107 3011 111
rect 3015 107 3017 111
rect 3021 107 3023 111
rect 3027 107 3029 111
rect 3033 107 3035 111
rect 3039 107 3383 111
rect 3387 107 3389 111
rect 3393 107 3395 111
rect 3399 107 3401 111
rect 3405 107 3407 111
rect 3411 107 3413 111
rect 3417 107 3419 111
rect 3423 107 3473 111
rect 3477 107 3479 111
rect 3483 107 3485 111
rect 3489 107 3491 111
rect 3495 107 3497 111
rect 3501 107 3503 111
rect 3507 107 3509 111
rect 3513 107 3857 111
rect 3861 107 3863 111
rect 3867 107 3869 111
rect 3873 107 3875 111
rect 3879 107 3881 111
rect 3885 107 3887 111
rect 3891 107 3893 111
rect 3897 107 3947 111
rect 3951 107 3953 111
rect 3957 107 3959 111
rect 3963 107 3965 111
rect 3969 107 3971 111
rect 3975 107 3977 111
rect 3981 107 3983 111
rect 3987 107 4331 111
rect 4335 107 4337 111
rect 4341 107 4343 111
rect 4347 107 4349 111
rect 4353 107 4355 111
rect 4359 107 4361 111
rect 4365 107 4367 111
rect 4371 107 4421 111
rect 4425 107 4427 111
rect 4431 107 4433 111
rect 4437 107 4439 111
rect 4443 107 4445 111
rect 4449 107 4451 111
rect 4455 107 4457 111
rect 4461 107 4633 111
rect 367 106 4633 107
rect 411 101 4589 102
rect 411 99 495 101
rect 411 65 413 99
rect 487 92 495 99
rect 499 92 501 101
rect 505 92 507 101
rect 511 92 513 101
rect 517 92 519 101
rect 523 92 525 101
rect 529 92 531 101
rect 535 92 673 101
rect 677 92 679 101
rect 683 92 685 101
rect 689 92 691 101
rect 695 92 697 101
rect 701 92 703 101
rect 707 92 709 101
rect 713 92 969 101
rect 973 92 975 101
rect 979 92 981 101
rect 985 92 987 101
rect 991 92 993 101
rect 997 92 999 101
rect 1003 92 1005 101
rect 1009 92 1147 101
rect 1151 92 1153 101
rect 1157 92 1159 101
rect 1163 92 1165 101
rect 1169 92 1171 101
rect 1175 92 1177 101
rect 1181 92 1183 101
rect 1187 92 1443 101
rect 1447 92 1449 101
rect 1453 92 1455 101
rect 1459 92 1461 101
rect 1465 92 1467 101
rect 1471 92 1473 101
rect 1477 92 1479 101
rect 1483 92 1621 101
rect 1625 92 1627 101
rect 1631 92 1633 101
rect 1637 92 1639 101
rect 1643 92 1645 101
rect 1649 92 1651 101
rect 1655 92 1657 101
rect 1661 92 1917 101
rect 1921 92 1923 101
rect 1927 92 1929 101
rect 1933 92 1935 101
rect 1939 92 1941 101
rect 1945 92 1947 101
rect 1951 92 1953 101
rect 1957 92 2095 101
rect 2099 92 2101 101
rect 2105 92 2107 101
rect 2111 92 2113 101
rect 2117 92 2119 101
rect 2123 92 2125 101
rect 2129 92 2131 101
rect 2135 92 2391 101
rect 2395 92 2397 101
rect 2401 92 2403 101
rect 2407 92 2409 101
rect 2413 92 2415 101
rect 2419 92 2421 101
rect 2425 92 2427 101
rect 2431 92 2569 101
rect 2573 92 2575 101
rect 2579 92 2581 101
rect 2585 92 2587 101
rect 2591 92 2593 101
rect 2597 92 2599 101
rect 2603 92 2605 101
rect 2609 92 2865 101
rect 2869 92 2871 101
rect 2875 92 2877 101
rect 2881 92 2883 101
rect 2887 92 2889 101
rect 2893 92 2895 101
rect 2899 92 2901 101
rect 2905 92 3043 101
rect 3047 92 3049 101
rect 3053 92 3055 101
rect 3059 92 3061 101
rect 3065 92 3067 101
rect 3071 92 3073 101
rect 3077 92 3079 101
rect 3083 92 3339 101
rect 3343 92 3345 101
rect 3349 92 3351 101
rect 3355 92 3357 101
rect 3361 92 3363 101
rect 3367 92 3369 101
rect 3373 92 3375 101
rect 3379 92 3517 101
rect 3521 92 3523 101
rect 3527 92 3529 101
rect 3533 92 3535 101
rect 3539 92 3541 101
rect 3545 92 3547 101
rect 3551 92 3553 101
rect 3557 92 3813 101
rect 3817 92 3819 101
rect 3823 92 3825 101
rect 3829 92 3831 101
rect 3835 92 3837 101
rect 3841 92 3843 101
rect 3847 92 3849 101
rect 3853 92 3991 101
rect 3995 92 3997 101
rect 4001 92 4003 101
rect 4007 92 4009 101
rect 4013 92 4015 101
rect 4019 92 4021 101
rect 4025 92 4027 101
rect 4031 92 4287 101
rect 4291 92 4293 101
rect 4297 92 4299 101
rect 4303 92 4305 101
rect 4309 92 4311 101
rect 4315 92 4317 101
rect 4321 92 4323 101
rect 4327 92 4465 101
rect 4469 92 4471 101
rect 4475 92 4477 101
rect 4481 92 4483 101
rect 4487 92 4489 101
rect 4493 92 4495 101
rect 4499 92 4501 101
rect 4505 92 4589 101
rect 487 90 4589 92
rect 487 86 495 90
rect 499 86 501 90
rect 505 86 507 90
rect 511 86 513 90
rect 517 86 519 90
rect 523 86 525 90
rect 529 86 531 90
rect 535 86 673 90
rect 677 86 679 90
rect 683 86 685 90
rect 689 86 691 90
rect 695 86 697 90
rect 701 86 703 90
rect 707 86 709 90
rect 713 86 969 90
rect 973 86 975 90
rect 979 86 981 90
rect 985 86 987 90
rect 991 86 993 90
rect 997 86 999 90
rect 1003 86 1005 90
rect 1009 86 1147 90
rect 1151 86 1153 90
rect 1157 86 1159 90
rect 1163 86 1165 90
rect 1169 86 1171 90
rect 1175 86 1177 90
rect 1181 86 1183 90
rect 1187 86 1443 90
rect 1447 86 1449 90
rect 1453 86 1455 90
rect 1459 86 1461 90
rect 1465 86 1467 90
rect 1471 86 1473 90
rect 1477 86 1479 90
rect 1483 86 1621 90
rect 1625 86 1627 90
rect 1631 86 1633 90
rect 1637 86 1639 90
rect 1643 86 1645 90
rect 1649 86 1651 90
rect 1655 86 1657 90
rect 1661 86 1917 90
rect 1921 86 1923 90
rect 1927 86 1929 90
rect 1933 86 1935 90
rect 1939 86 1941 90
rect 1945 86 1947 90
rect 1951 86 1953 90
rect 1957 86 2095 90
rect 2099 86 2101 90
rect 2105 86 2107 90
rect 2111 86 2113 90
rect 2117 86 2119 90
rect 2123 86 2125 90
rect 2129 86 2131 90
rect 2135 86 2391 90
rect 2395 86 2397 90
rect 2401 86 2403 90
rect 2407 86 2409 90
rect 2413 86 2415 90
rect 2419 86 2421 90
rect 2425 86 2427 90
rect 2431 86 2569 90
rect 2573 86 2575 90
rect 2579 86 2581 90
rect 2585 86 2587 90
rect 2591 86 2593 90
rect 2597 86 2599 90
rect 2603 86 2605 90
rect 2609 86 2865 90
rect 2869 86 2871 90
rect 2875 86 2877 90
rect 2881 86 2883 90
rect 2887 86 2889 90
rect 2893 86 2895 90
rect 2899 86 2901 90
rect 2905 86 3043 90
rect 3047 86 3049 90
rect 3053 86 3055 90
rect 3059 86 3061 90
rect 3065 86 3067 90
rect 3071 86 3073 90
rect 3077 86 3079 90
rect 3083 86 3339 90
rect 3343 86 3345 90
rect 3349 86 3351 90
rect 3355 86 3357 90
rect 3361 86 3363 90
rect 3367 86 3369 90
rect 3373 86 3375 90
rect 3379 86 3517 90
rect 3521 86 3523 90
rect 3527 86 3529 90
rect 3533 86 3535 90
rect 3539 86 3541 90
rect 3545 86 3547 90
rect 3551 86 3553 90
rect 3557 86 3813 90
rect 3817 86 3819 90
rect 3823 86 3825 90
rect 3829 86 3831 90
rect 3835 86 3837 90
rect 3841 86 3843 90
rect 3847 86 3849 90
rect 3853 86 3991 90
rect 3995 86 3997 90
rect 4001 86 4003 90
rect 4007 86 4009 90
rect 4013 86 4015 90
rect 4019 86 4021 90
rect 4025 86 4027 90
rect 4031 86 4287 90
rect 4291 86 4293 90
rect 4297 86 4299 90
rect 4303 86 4305 90
rect 4309 86 4311 90
rect 4315 86 4317 90
rect 4321 86 4323 90
rect 4327 86 4465 90
rect 4469 86 4471 90
rect 4475 86 4477 90
rect 4481 86 4483 90
rect 4487 86 4489 90
rect 4493 86 4495 90
rect 4499 86 4501 90
rect 4505 86 4589 90
rect 487 84 4589 86
rect 487 80 495 84
rect 499 80 501 84
rect 505 80 507 84
rect 511 80 513 84
rect 517 80 519 84
rect 523 80 525 84
rect 529 80 531 84
rect 535 80 673 84
rect 677 80 679 84
rect 683 80 685 84
rect 689 80 691 84
rect 695 80 697 84
rect 701 80 703 84
rect 707 80 709 84
rect 713 80 969 84
rect 973 80 975 84
rect 979 80 981 84
rect 985 80 987 84
rect 991 80 993 84
rect 997 80 999 84
rect 1003 80 1005 84
rect 1009 80 1147 84
rect 1151 80 1153 84
rect 1157 80 1159 84
rect 1163 80 1165 84
rect 1169 80 1171 84
rect 1175 80 1177 84
rect 1181 80 1183 84
rect 1187 80 1443 84
rect 1447 80 1449 84
rect 1453 80 1455 84
rect 1459 80 1461 84
rect 1465 80 1467 84
rect 1471 80 1473 84
rect 1477 80 1479 84
rect 1483 80 1621 84
rect 1625 80 1627 84
rect 1631 80 1633 84
rect 1637 80 1639 84
rect 1643 80 1645 84
rect 1649 80 1651 84
rect 1655 80 1657 84
rect 1661 80 1917 84
rect 1921 80 1923 84
rect 1927 80 1929 84
rect 1933 80 1935 84
rect 1939 80 1941 84
rect 1945 80 1947 84
rect 1951 80 1953 84
rect 1957 80 2095 84
rect 2099 80 2101 84
rect 2105 80 2107 84
rect 2111 80 2113 84
rect 2117 80 2119 84
rect 2123 80 2125 84
rect 2129 80 2131 84
rect 2135 80 2391 84
rect 2395 80 2397 84
rect 2401 80 2403 84
rect 2407 80 2409 84
rect 2413 80 2415 84
rect 2419 80 2421 84
rect 2425 80 2427 84
rect 2431 80 2569 84
rect 2573 80 2575 84
rect 2579 80 2581 84
rect 2585 80 2587 84
rect 2591 80 2593 84
rect 2597 80 2599 84
rect 2603 80 2605 84
rect 2609 80 2865 84
rect 2869 80 2871 84
rect 2875 80 2877 84
rect 2881 80 2883 84
rect 2887 80 2889 84
rect 2893 80 2895 84
rect 2899 80 2901 84
rect 2905 80 3043 84
rect 3047 80 3049 84
rect 3053 80 3055 84
rect 3059 80 3061 84
rect 3065 80 3067 84
rect 3071 80 3073 84
rect 3077 80 3079 84
rect 3083 80 3339 84
rect 3343 80 3345 84
rect 3349 80 3351 84
rect 3355 80 3357 84
rect 3361 80 3363 84
rect 3367 80 3369 84
rect 3373 80 3375 84
rect 3379 80 3517 84
rect 3521 80 3523 84
rect 3527 80 3529 84
rect 3533 80 3535 84
rect 3539 80 3541 84
rect 3545 80 3547 84
rect 3551 80 3553 84
rect 3557 80 3813 84
rect 3817 80 3819 84
rect 3823 80 3825 84
rect 3829 80 3831 84
rect 3835 80 3837 84
rect 3841 80 3843 84
rect 3847 80 3849 84
rect 3853 80 3991 84
rect 3995 80 3997 84
rect 4001 80 4003 84
rect 4007 80 4009 84
rect 4013 80 4015 84
rect 4019 80 4021 84
rect 4025 80 4027 84
rect 4031 80 4287 84
rect 4291 80 4293 84
rect 4297 80 4299 84
rect 4303 80 4305 84
rect 4309 80 4311 84
rect 4315 80 4317 84
rect 4321 80 4323 84
rect 4327 80 4465 84
rect 4469 80 4471 84
rect 4475 80 4477 84
rect 4481 80 4483 84
rect 4487 80 4489 84
rect 4493 80 4495 84
rect 4499 80 4501 84
rect 4505 80 4589 84
rect 487 78 4589 80
rect 487 74 495 78
rect 499 74 501 78
rect 505 74 507 78
rect 511 74 513 78
rect 517 74 519 78
rect 523 74 525 78
rect 529 74 531 78
rect 535 74 673 78
rect 677 74 679 78
rect 683 74 685 78
rect 689 74 691 78
rect 695 74 697 78
rect 701 74 703 78
rect 707 74 709 78
rect 713 74 969 78
rect 973 74 975 78
rect 979 74 981 78
rect 985 74 987 78
rect 991 74 993 78
rect 997 74 999 78
rect 1003 74 1005 78
rect 1009 74 1147 78
rect 1151 74 1153 78
rect 1157 74 1159 78
rect 1163 74 1165 78
rect 1169 74 1171 78
rect 1175 74 1177 78
rect 1181 74 1183 78
rect 1187 74 1443 78
rect 1447 74 1449 78
rect 1453 74 1455 78
rect 1459 74 1461 78
rect 1465 74 1467 78
rect 1471 74 1473 78
rect 1477 74 1479 78
rect 1483 74 1621 78
rect 1625 74 1627 78
rect 1631 74 1633 78
rect 1637 74 1639 78
rect 1643 74 1645 78
rect 1649 74 1651 78
rect 1655 74 1657 78
rect 1661 74 1917 78
rect 1921 74 1923 78
rect 1927 74 1929 78
rect 1933 74 1935 78
rect 1939 74 1941 78
rect 1945 74 1947 78
rect 1951 74 1953 78
rect 1957 74 2095 78
rect 2099 74 2101 78
rect 2105 74 2107 78
rect 2111 74 2113 78
rect 2117 74 2119 78
rect 2123 74 2125 78
rect 2129 74 2131 78
rect 2135 74 2391 78
rect 2395 74 2397 78
rect 2401 74 2403 78
rect 2407 74 2409 78
rect 2413 74 2415 78
rect 2419 74 2421 78
rect 2425 74 2427 78
rect 2431 74 2569 78
rect 2573 74 2575 78
rect 2579 74 2581 78
rect 2585 74 2587 78
rect 2591 74 2593 78
rect 2597 74 2599 78
rect 2603 74 2605 78
rect 2609 74 2865 78
rect 2869 74 2871 78
rect 2875 74 2877 78
rect 2881 74 2883 78
rect 2887 74 2889 78
rect 2893 74 2895 78
rect 2899 74 2901 78
rect 2905 74 3043 78
rect 3047 74 3049 78
rect 3053 74 3055 78
rect 3059 74 3061 78
rect 3065 74 3067 78
rect 3071 74 3073 78
rect 3077 74 3079 78
rect 3083 74 3339 78
rect 3343 74 3345 78
rect 3349 74 3351 78
rect 3355 74 3357 78
rect 3361 74 3363 78
rect 3367 74 3369 78
rect 3373 74 3375 78
rect 3379 74 3517 78
rect 3521 74 3523 78
rect 3527 74 3529 78
rect 3533 74 3535 78
rect 3539 74 3541 78
rect 3545 74 3547 78
rect 3551 74 3553 78
rect 3557 74 3813 78
rect 3817 74 3819 78
rect 3823 74 3825 78
rect 3829 74 3831 78
rect 3835 74 3837 78
rect 3841 74 3843 78
rect 3847 74 3849 78
rect 3853 74 3991 78
rect 3995 74 3997 78
rect 4001 74 4003 78
rect 4007 74 4009 78
rect 4013 74 4015 78
rect 4019 74 4021 78
rect 4025 74 4027 78
rect 4031 74 4287 78
rect 4291 74 4293 78
rect 4297 74 4299 78
rect 4303 74 4305 78
rect 4309 74 4311 78
rect 4315 74 4317 78
rect 4321 74 4323 78
rect 4327 74 4465 78
rect 4469 74 4471 78
rect 4475 74 4477 78
rect 4481 74 4483 78
rect 4487 74 4489 78
rect 4493 74 4495 78
rect 4499 74 4501 78
rect 4505 74 4589 78
rect 487 72 4589 74
rect 487 65 495 72
rect 411 63 495 65
rect 499 63 501 72
rect 505 63 507 72
rect 511 63 513 72
rect 517 63 519 72
rect 523 63 525 72
rect 529 63 531 72
rect 535 63 673 72
rect 677 63 679 72
rect 683 63 685 72
rect 689 63 691 72
rect 695 63 697 72
rect 701 63 703 72
rect 707 63 709 72
rect 713 63 969 72
rect 973 63 975 72
rect 979 63 981 72
rect 985 63 987 72
rect 991 63 993 72
rect 997 63 999 72
rect 1003 63 1005 72
rect 1009 63 1147 72
rect 1151 63 1153 72
rect 1157 63 1159 72
rect 1163 63 1165 72
rect 1169 63 1171 72
rect 1175 63 1177 72
rect 1181 63 1183 72
rect 1187 63 1443 72
rect 1447 63 1449 72
rect 1453 63 1455 72
rect 1459 63 1461 72
rect 1465 63 1467 72
rect 1471 63 1473 72
rect 1477 63 1479 72
rect 1483 63 1621 72
rect 1625 63 1627 72
rect 1631 63 1633 72
rect 1637 63 1639 72
rect 1643 63 1645 72
rect 1649 63 1651 72
rect 1655 63 1657 72
rect 1661 63 1917 72
rect 1921 63 1923 72
rect 1927 63 1929 72
rect 1933 63 1935 72
rect 1939 63 1941 72
rect 1945 63 1947 72
rect 1951 63 1953 72
rect 1957 63 2095 72
rect 2099 63 2101 72
rect 2105 63 2107 72
rect 2111 63 2113 72
rect 2117 63 2119 72
rect 2123 63 2125 72
rect 2129 63 2131 72
rect 2135 63 2391 72
rect 2395 63 2397 72
rect 2401 63 2403 72
rect 2407 63 2409 72
rect 2413 63 2415 72
rect 2419 63 2421 72
rect 2425 63 2427 72
rect 2431 63 2569 72
rect 2573 63 2575 72
rect 2579 63 2581 72
rect 2585 63 2587 72
rect 2591 63 2593 72
rect 2597 63 2599 72
rect 2603 63 2605 72
rect 2609 63 2865 72
rect 2869 63 2871 72
rect 2875 63 2877 72
rect 2881 63 2883 72
rect 2887 63 2889 72
rect 2893 63 2895 72
rect 2899 63 2901 72
rect 2905 63 3043 72
rect 3047 63 3049 72
rect 3053 63 3055 72
rect 3059 63 3061 72
rect 3065 63 3067 72
rect 3071 63 3073 72
rect 3077 63 3079 72
rect 3083 63 3339 72
rect 3343 63 3345 72
rect 3349 63 3351 72
rect 3355 63 3357 72
rect 3361 63 3363 72
rect 3367 63 3369 72
rect 3373 63 3375 72
rect 3379 63 3517 72
rect 3521 63 3523 72
rect 3527 63 3529 72
rect 3533 63 3535 72
rect 3539 63 3541 72
rect 3545 63 3547 72
rect 3551 63 3553 72
rect 3557 63 3813 72
rect 3817 63 3819 72
rect 3823 63 3825 72
rect 3829 63 3831 72
rect 3835 63 3837 72
rect 3841 63 3843 72
rect 3847 63 3849 72
rect 3853 63 3991 72
rect 3995 63 3997 72
rect 4001 63 4003 72
rect 4007 63 4009 72
rect 4013 63 4015 72
rect 4019 63 4021 72
rect 4025 63 4027 72
rect 4031 63 4287 72
rect 4291 63 4293 72
rect 4297 63 4299 72
rect 4303 63 4305 72
rect 4309 63 4311 72
rect 4315 63 4317 72
rect 4321 63 4323 72
rect 4327 63 4465 72
rect 4469 63 4471 72
rect 4475 63 4477 72
rect 4481 63 4483 72
rect 4487 63 4489 72
rect 4493 63 4495 72
rect 4499 63 4501 72
rect 4505 63 4589 72
rect 411 62 4589 63
rect 455 57 4545 58
rect 455 53 578 57
rect 582 53 588 57
rect 592 53 616 57
rect 620 53 626 57
rect 630 53 1052 57
rect 1056 53 1062 57
rect 1066 53 1090 57
rect 1094 53 1100 57
rect 1104 53 1526 57
rect 1530 53 1536 57
rect 1540 53 1564 57
rect 1568 53 1574 57
rect 1578 53 2000 57
rect 2004 53 2010 57
rect 2014 53 2038 57
rect 2042 53 2048 57
rect 2052 53 2474 57
rect 2478 53 2484 57
rect 2488 53 2512 57
rect 2516 53 2522 57
rect 2526 53 2948 57
rect 2952 53 2958 57
rect 2962 53 2986 57
rect 2990 53 2996 57
rect 3000 53 3422 57
rect 3426 53 3432 57
rect 3436 53 3460 57
rect 3464 53 3470 57
rect 3474 53 3896 57
rect 3900 53 3906 57
rect 3910 53 3934 57
rect 3938 53 3944 57
rect 3948 53 4370 57
rect 4374 53 4380 57
rect 4384 53 4408 57
rect 4412 53 4418 57
rect 4422 53 4470 57
rect 4544 53 4545 57
rect 455 52 4545 53
rect 465 47 1013 48
rect 465 43 539 47
rect 543 43 545 47
rect 549 43 551 47
rect 555 43 557 47
rect 561 43 563 47
rect 567 43 569 47
rect 573 43 575 47
rect 579 43 629 47
rect 633 43 635 47
rect 639 43 641 47
rect 645 43 647 47
rect 651 43 653 47
rect 657 43 659 47
rect 663 43 665 47
rect 669 44 1013 47
rect 1017 44 1019 48
rect 1023 44 1025 48
rect 1029 44 1031 48
rect 1035 44 1037 48
rect 1041 44 1043 48
rect 1047 44 1049 48
rect 1053 44 1103 48
rect 1107 44 1109 48
rect 1113 44 1115 48
rect 1119 44 1121 48
rect 1125 44 1127 48
rect 1131 44 1133 48
rect 1137 44 1139 48
rect 1143 44 1487 48
rect 1491 44 1493 48
rect 1497 44 1499 48
rect 1503 44 1505 48
rect 1509 44 1511 48
rect 1515 44 1517 48
rect 1521 44 1523 48
rect 1527 44 1577 48
rect 1581 44 1583 48
rect 1587 44 1589 48
rect 1593 44 1595 48
rect 1599 44 1601 48
rect 1605 44 1607 48
rect 1611 44 1613 48
rect 1617 44 1961 48
rect 1965 44 1967 48
rect 1971 44 1973 48
rect 1977 44 1979 48
rect 1983 44 1985 48
rect 1989 44 1991 48
rect 1995 44 1997 48
rect 2001 44 2051 48
rect 2055 44 2057 48
rect 2061 44 2063 48
rect 2067 44 2069 48
rect 2073 44 2075 48
rect 2079 44 2081 48
rect 2085 44 2087 48
rect 2091 44 2435 48
rect 2439 44 2441 48
rect 2445 44 2447 48
rect 2451 44 2453 48
rect 2457 44 2459 48
rect 2463 44 2465 48
rect 2469 44 2471 48
rect 2475 44 2525 48
rect 2529 44 2531 48
rect 2535 44 2537 48
rect 2541 44 2543 48
rect 2547 44 2549 48
rect 2553 44 2555 48
rect 2559 44 2561 48
rect 2565 44 2909 48
rect 2913 44 2915 48
rect 2919 44 2921 48
rect 2925 44 2927 48
rect 2931 44 2933 48
rect 2937 44 2939 48
rect 2943 44 2945 48
rect 2949 44 2999 48
rect 3003 44 3005 48
rect 3009 44 3011 48
rect 3015 44 3017 48
rect 3021 44 3023 48
rect 3027 44 3029 48
rect 3033 44 3035 48
rect 3039 44 3383 48
rect 3387 44 3389 48
rect 3393 44 3395 48
rect 3399 44 3401 48
rect 3405 44 3407 48
rect 3411 44 3413 48
rect 3417 44 3419 48
rect 3423 44 3473 48
rect 3477 44 3479 48
rect 3483 44 3485 48
rect 3489 44 3491 48
rect 3495 44 3497 48
rect 3501 44 3503 48
rect 3507 44 3509 48
rect 3513 44 3857 48
rect 3861 44 3863 48
rect 3867 44 3869 48
rect 3873 44 3875 48
rect 3879 44 3881 48
rect 3885 44 3887 48
rect 3891 44 3893 48
rect 3897 44 3947 48
rect 3951 44 3953 48
rect 3957 44 3959 48
rect 3963 44 3965 48
rect 3969 44 3971 48
rect 3975 44 3977 48
rect 3981 44 3983 48
rect 3987 44 4331 48
rect 4335 44 4337 48
rect 4341 44 4343 48
rect 4347 44 4349 48
rect 4353 44 4355 48
rect 4359 44 4361 48
rect 4365 44 4367 48
rect 4371 44 4421 48
rect 4425 44 4427 48
rect 4431 44 4433 48
rect 4437 44 4439 48
rect 4443 44 4445 48
rect 4449 44 4451 48
rect 4455 44 4457 48
rect 4461 44 4535 48
rect 669 43 4535 44
rect 465 36 4535 43
rect 465 32 539 36
rect 543 32 545 36
rect 549 32 551 36
rect 555 32 557 36
rect 561 32 563 36
rect 567 32 569 36
rect 573 32 575 36
rect 579 32 629 36
rect 633 32 635 36
rect 639 32 641 36
rect 645 32 647 36
rect 651 32 653 36
rect 657 32 659 36
rect 663 32 665 36
rect 669 32 1013 36
rect 1017 32 1019 36
rect 1023 32 1025 36
rect 1029 32 1031 36
rect 1035 32 1037 36
rect 1041 32 1043 36
rect 1047 32 1049 36
rect 1053 32 1103 36
rect 1107 32 1109 36
rect 1113 32 1115 36
rect 1119 32 1121 36
rect 1125 32 1127 36
rect 1131 32 1133 36
rect 1137 32 1139 36
rect 1143 32 1487 36
rect 1491 32 1493 36
rect 1497 32 1499 36
rect 1503 32 1505 36
rect 1509 32 1511 36
rect 1515 32 1517 36
rect 1521 32 1523 36
rect 1527 32 1577 36
rect 1581 32 1583 36
rect 1587 32 1589 36
rect 1593 32 1595 36
rect 1599 32 1601 36
rect 1605 32 1607 36
rect 1611 32 1613 36
rect 1617 32 1961 36
rect 1965 32 1967 36
rect 1971 32 1973 36
rect 1977 32 1979 36
rect 1983 32 1985 36
rect 1989 32 1991 36
rect 1995 32 1997 36
rect 2001 32 2051 36
rect 2055 32 2057 36
rect 2061 32 2063 36
rect 2067 32 2069 36
rect 2073 32 2075 36
rect 2079 32 2081 36
rect 2085 32 2087 36
rect 2091 32 2435 36
rect 2439 32 2441 36
rect 2445 32 2447 36
rect 2451 32 2453 36
rect 2457 32 2459 36
rect 2463 32 2465 36
rect 2469 32 2471 36
rect 2475 32 2525 36
rect 2529 32 2531 36
rect 2535 32 2537 36
rect 2541 32 2543 36
rect 2547 32 2549 36
rect 2553 32 2555 36
rect 2559 32 2561 36
rect 2565 32 2909 36
rect 2913 32 2915 36
rect 2919 32 2921 36
rect 2925 32 2927 36
rect 2931 32 2933 36
rect 2937 32 2939 36
rect 2943 32 2945 36
rect 2949 32 2999 36
rect 3003 32 3005 36
rect 3009 32 3011 36
rect 3015 32 3017 36
rect 3021 32 3023 36
rect 3027 32 3029 36
rect 3033 32 3035 36
rect 3039 32 3383 36
rect 3387 32 3389 36
rect 3393 32 3395 36
rect 3399 32 3401 36
rect 3405 32 3407 36
rect 3411 32 3413 36
rect 3417 32 3419 36
rect 3423 32 3473 36
rect 3477 32 3479 36
rect 3483 32 3485 36
rect 3489 32 3491 36
rect 3495 32 3497 36
rect 3501 32 3503 36
rect 3507 32 3509 36
rect 3513 32 3857 36
rect 3861 32 3863 36
rect 3867 32 3869 36
rect 3873 32 3875 36
rect 3879 32 3881 36
rect 3885 32 3887 36
rect 3891 32 3893 36
rect 3897 32 3947 36
rect 3951 32 3953 36
rect 3957 32 3959 36
rect 3963 32 3965 36
rect 3969 32 3971 36
rect 3975 32 3977 36
rect 3981 32 3983 36
rect 3987 32 4331 36
rect 4335 32 4337 36
rect 4341 32 4343 36
rect 4347 32 4349 36
rect 4353 32 4355 36
rect 4359 32 4361 36
rect 4365 32 4367 36
rect 4371 32 4421 36
rect 4425 32 4427 36
rect 4431 32 4433 36
rect 4437 32 4439 36
rect 4443 32 4445 36
rect 4449 32 4451 36
rect 4455 32 4457 36
rect 4461 32 4535 36
rect 465 30 4535 32
rect 465 26 539 30
rect 543 26 545 30
rect 549 26 551 30
rect 555 26 557 30
rect 561 26 563 30
rect 567 26 569 30
rect 573 26 575 30
rect 579 26 629 30
rect 633 26 635 30
rect 639 26 641 30
rect 645 26 647 30
rect 651 26 653 30
rect 657 26 659 30
rect 663 26 665 30
rect 669 26 1013 30
rect 1017 26 1019 30
rect 1023 26 1025 30
rect 1029 26 1031 30
rect 1035 26 1037 30
rect 1041 26 1043 30
rect 1047 26 1049 30
rect 1053 26 1103 30
rect 1107 26 1109 30
rect 1113 26 1115 30
rect 1119 26 1121 30
rect 1125 26 1127 30
rect 1131 26 1133 30
rect 1137 26 1139 30
rect 1143 26 1487 30
rect 1491 26 1493 30
rect 1497 26 1499 30
rect 1503 26 1505 30
rect 1509 26 1511 30
rect 1515 26 1517 30
rect 1521 26 1523 30
rect 1527 26 1577 30
rect 1581 26 1583 30
rect 1587 26 1589 30
rect 1593 26 1595 30
rect 1599 26 1601 30
rect 1605 26 1607 30
rect 1611 26 1613 30
rect 1617 26 1961 30
rect 1965 26 1967 30
rect 1971 26 1973 30
rect 1977 26 1979 30
rect 1983 26 1985 30
rect 1989 26 1991 30
rect 1995 26 1997 30
rect 2001 26 2051 30
rect 2055 26 2057 30
rect 2061 26 2063 30
rect 2067 26 2069 30
rect 2073 26 2075 30
rect 2079 26 2081 30
rect 2085 26 2087 30
rect 2091 26 2435 30
rect 2439 26 2441 30
rect 2445 26 2447 30
rect 2451 26 2453 30
rect 2457 26 2459 30
rect 2463 26 2465 30
rect 2469 26 2471 30
rect 2475 26 2525 30
rect 2529 26 2531 30
rect 2535 26 2537 30
rect 2541 26 2543 30
rect 2547 26 2549 30
rect 2553 26 2555 30
rect 2559 26 2561 30
rect 2565 26 2909 30
rect 2913 26 2915 30
rect 2919 26 2921 30
rect 2925 26 2927 30
rect 2931 26 2933 30
rect 2937 26 2939 30
rect 2943 26 2945 30
rect 2949 26 2999 30
rect 3003 26 3005 30
rect 3009 26 3011 30
rect 3015 26 3017 30
rect 3021 26 3023 30
rect 3027 26 3029 30
rect 3033 26 3035 30
rect 3039 26 3383 30
rect 3387 26 3389 30
rect 3393 26 3395 30
rect 3399 26 3401 30
rect 3405 26 3407 30
rect 3411 26 3413 30
rect 3417 26 3419 30
rect 3423 26 3473 30
rect 3477 26 3479 30
rect 3483 26 3485 30
rect 3489 26 3491 30
rect 3495 26 3497 30
rect 3501 26 3503 30
rect 3507 26 3509 30
rect 3513 26 3857 30
rect 3861 26 3863 30
rect 3867 26 3869 30
rect 3873 26 3875 30
rect 3879 26 3881 30
rect 3885 26 3887 30
rect 3891 26 3893 30
rect 3897 26 3947 30
rect 3951 26 3953 30
rect 3957 26 3959 30
rect 3963 26 3965 30
rect 3969 26 3971 30
rect 3975 26 3977 30
rect 3981 26 3983 30
rect 3987 26 4331 30
rect 4335 26 4337 30
rect 4341 26 4343 30
rect 4347 26 4349 30
rect 4353 26 4355 30
rect 4359 26 4361 30
rect 4365 26 4367 30
rect 4371 26 4421 30
rect 4425 26 4427 30
rect 4431 26 4433 30
rect 4437 26 4439 30
rect 4443 26 4445 30
rect 4449 26 4451 30
rect 4455 26 4457 30
rect 4461 26 4535 30
rect 465 18 4535 26
rect 465 14 539 18
rect 543 14 545 18
rect 549 14 551 18
rect 555 14 557 18
rect 561 14 563 18
rect 567 14 569 18
rect 573 14 575 18
rect 579 14 629 18
rect 633 14 635 18
rect 639 14 641 18
rect 645 14 647 18
rect 651 14 653 18
rect 657 14 659 18
rect 663 14 1019 18
rect 1023 14 1025 18
rect 1029 14 1031 18
rect 1035 14 1037 18
rect 1041 14 1043 18
rect 1047 14 1049 18
rect 1053 14 1103 18
rect 1107 14 1109 18
rect 1113 14 1115 18
rect 1119 14 1121 18
rect 1125 14 1127 18
rect 1131 14 1133 18
rect 1137 14 1493 18
rect 1497 14 1499 18
rect 1503 14 1505 18
rect 1509 14 1511 18
rect 1515 14 1517 18
rect 1521 14 1523 18
rect 1527 14 1577 18
rect 1581 14 1583 18
rect 1587 14 1589 18
rect 1593 14 1595 18
rect 1599 14 1601 18
rect 1605 14 1607 18
rect 1611 14 1967 18
rect 1971 14 1973 18
rect 1977 14 1979 18
rect 1983 14 1985 18
rect 1989 14 1991 18
rect 1995 14 1997 18
rect 2001 14 2051 18
rect 2055 14 2057 18
rect 2061 14 2063 18
rect 2067 14 2069 18
rect 2073 14 2075 18
rect 2079 14 2081 18
rect 2085 14 2441 18
rect 2445 14 2447 18
rect 2451 14 2453 18
rect 2457 14 2459 18
rect 2463 14 2465 18
rect 2469 14 2471 18
rect 2475 14 2525 18
rect 2529 14 2531 18
rect 2535 14 2537 18
rect 2541 14 2543 18
rect 2547 14 2549 18
rect 2553 14 2555 18
rect 2559 14 2915 18
rect 2919 14 2921 18
rect 2925 14 2927 18
rect 2931 14 2933 18
rect 2937 14 2939 18
rect 2943 14 2945 18
rect 2949 14 2999 18
rect 3003 14 3005 18
rect 3009 14 3011 18
rect 3015 14 3017 18
rect 3021 14 3023 18
rect 3027 14 3029 18
rect 3033 14 3389 18
rect 3393 14 3395 18
rect 3399 14 3401 18
rect 3405 14 3407 18
rect 3411 14 3413 18
rect 3417 14 3419 18
rect 3423 14 3473 18
rect 3477 14 3479 18
rect 3483 14 3485 18
rect 3489 14 3491 18
rect 3495 14 3497 18
rect 3501 14 3503 18
rect 3507 14 3863 18
rect 3867 14 3869 18
rect 3873 14 3875 18
rect 3879 14 3881 18
rect 3885 14 3887 18
rect 3891 14 3893 18
rect 3897 14 3947 18
rect 3951 14 3953 18
rect 3957 14 3959 18
rect 3963 14 3965 18
rect 3969 14 3971 18
rect 3975 14 3977 18
rect 3981 14 4337 18
rect 4341 14 4343 18
rect 4347 14 4349 18
rect 4353 14 4355 18
rect 4359 14 4361 18
rect 4365 14 4367 18
rect 4371 14 4421 18
rect 4425 14 4427 18
rect 4431 14 4433 18
rect 4437 14 4439 18
rect 4443 14 4445 18
rect 4449 14 4451 18
rect 4455 14 4457 18
rect 4461 14 4535 18
rect 465 8 4535 14
rect 539 4 579 8
rect 629 4 669 8
rect 1013 4 1053 8
rect 1103 4 1143 8
rect 1487 4 1527 8
rect 1577 4 1617 8
rect 1961 4 2001 8
rect 2051 4 2091 8
rect 2435 4 2475 8
rect 2525 4 2565 8
rect 2909 4 2949 8
rect 2999 4 3039 8
rect 3383 4 3423 8
rect 3473 4 3513 8
rect 3857 4 3897 8
rect 3947 4 3987 8
rect 4331 4 4371 8
rect 4421 4 4461 8
rect 543 0 545 4
rect 549 0 551 4
rect 555 0 557 4
rect 561 0 563 4
rect 567 0 569 4
rect 573 0 575 4
rect 633 0 635 4
rect 639 0 641 4
rect 645 0 647 4
rect 651 0 653 4
rect 657 0 659 4
rect 663 0 665 4
rect 677 0 679 4
rect 683 0 685 4
rect 689 0 691 4
rect 695 0 697 4
rect 701 0 703 4
rect 707 0 709 4
rect 973 0 975 4
rect 979 0 981 4
rect 985 0 987 4
rect 991 0 993 4
rect 997 0 999 4
rect 1003 0 1005 4
rect 1017 0 1019 4
rect 1023 0 1025 4
rect 1029 0 1031 4
rect 1035 0 1037 4
rect 1041 0 1043 4
rect 1047 0 1049 4
rect 1107 0 1109 4
rect 1113 0 1115 4
rect 1119 0 1121 4
rect 1125 0 1127 4
rect 1131 0 1133 4
rect 1137 0 1139 4
rect 1151 0 1153 4
rect 1157 0 1159 4
rect 1163 0 1165 4
rect 1169 0 1171 4
rect 1175 0 1177 4
rect 1181 0 1183 4
rect 1447 0 1449 4
rect 1453 0 1455 4
rect 1459 0 1461 4
rect 1465 0 1467 4
rect 1471 0 1473 4
rect 1477 0 1479 4
rect 1491 0 1493 4
rect 1497 0 1499 4
rect 1503 0 1505 4
rect 1509 0 1511 4
rect 1515 0 1517 4
rect 1521 0 1523 4
rect 1581 0 1583 4
rect 1587 0 1589 4
rect 1593 0 1595 4
rect 1599 0 1601 4
rect 1605 0 1607 4
rect 1611 0 1613 4
rect 1625 0 1627 4
rect 1631 0 1633 4
rect 1637 0 1639 4
rect 1643 0 1645 4
rect 1649 0 1651 4
rect 1655 0 1657 4
rect 1921 0 1923 4
rect 1927 0 1929 4
rect 1933 0 1935 4
rect 1939 0 1941 4
rect 1945 0 1947 4
rect 1951 0 1953 4
rect 1965 0 1967 4
rect 1971 0 1973 4
rect 1977 0 1979 4
rect 1983 0 1985 4
rect 1989 0 1991 4
rect 1995 0 1997 4
rect 2055 0 2057 4
rect 2061 0 2063 4
rect 2067 0 2069 4
rect 2073 0 2075 4
rect 2079 0 2081 4
rect 2085 0 2087 4
rect 2099 0 2101 4
rect 2105 0 2107 4
rect 2111 0 2113 4
rect 2117 0 2119 4
rect 2123 0 2125 4
rect 2129 0 2131 4
rect 2395 0 2397 4
rect 2401 0 2403 4
rect 2407 0 2409 4
rect 2413 0 2415 4
rect 2419 0 2421 4
rect 2425 0 2427 4
rect 2439 0 2441 4
rect 2445 0 2447 4
rect 2451 0 2453 4
rect 2457 0 2459 4
rect 2463 0 2465 4
rect 2469 0 2471 4
rect 2529 0 2531 4
rect 2535 0 2537 4
rect 2541 0 2543 4
rect 2547 0 2549 4
rect 2553 0 2555 4
rect 2559 0 2561 4
rect 2573 0 2575 4
rect 2579 0 2581 4
rect 2585 0 2587 4
rect 2591 0 2593 4
rect 2597 0 2599 4
rect 2603 0 2605 4
rect 2869 0 2871 4
rect 2875 0 2877 4
rect 2881 0 2883 4
rect 2887 0 2889 4
rect 2893 0 2895 4
rect 2899 0 2901 4
rect 2913 0 2915 4
rect 2919 0 2921 4
rect 2925 0 2927 4
rect 2931 0 2933 4
rect 2937 0 2939 4
rect 2943 0 2945 4
rect 3003 0 3005 4
rect 3009 0 3011 4
rect 3015 0 3017 4
rect 3021 0 3023 4
rect 3027 0 3029 4
rect 3033 0 3035 4
rect 3047 0 3049 4
rect 3053 0 3055 4
rect 3059 0 3061 4
rect 3065 0 3067 4
rect 3071 0 3073 4
rect 3077 0 3079 4
rect 3343 0 3345 4
rect 3349 0 3351 4
rect 3355 0 3357 4
rect 3361 0 3363 4
rect 3367 0 3369 4
rect 3373 0 3375 4
rect 3387 0 3389 4
rect 3393 0 3395 4
rect 3399 0 3401 4
rect 3405 0 3407 4
rect 3411 0 3413 4
rect 3417 0 3419 4
rect 3477 0 3479 4
rect 3483 0 3485 4
rect 3489 0 3491 4
rect 3495 0 3497 4
rect 3501 0 3503 4
rect 3507 0 3509 4
rect 3521 0 3523 4
rect 3527 0 3529 4
rect 3533 0 3535 4
rect 3539 0 3541 4
rect 3545 0 3547 4
rect 3551 0 3553 4
rect 3817 0 3819 4
rect 3823 0 3825 4
rect 3829 0 3831 4
rect 3835 0 3837 4
rect 3841 0 3843 4
rect 3847 0 3849 4
rect 3861 0 3863 4
rect 3867 0 3869 4
rect 3873 0 3875 4
rect 3879 0 3881 4
rect 3885 0 3887 4
rect 3891 0 3893 4
rect 3951 0 3953 4
rect 3957 0 3959 4
rect 3963 0 3965 4
rect 3969 0 3971 4
rect 3975 0 3977 4
rect 3981 0 3983 4
rect 3995 0 3997 4
rect 4001 0 4003 4
rect 4007 0 4009 4
rect 4013 0 4015 4
rect 4019 0 4021 4
rect 4025 0 4027 4
rect 4291 0 4293 4
rect 4297 0 4299 4
rect 4303 0 4305 4
rect 4309 0 4311 4
rect 4315 0 4317 4
rect 4321 0 4323 4
rect 4335 0 4337 4
rect 4341 0 4343 4
rect 4347 0 4349 4
rect 4353 0 4355 4
rect 4359 0 4361 4
rect 4365 0 4367 4
rect 4425 0 4427 4
rect 4431 0 4433 4
rect 4437 0 4439 4
rect 4443 0 4445 4
rect 4449 0 4451 4
rect 4455 0 4457 4
<< m3contact >>
rect 4644 490 4653 499
rect 413 65 487 99
rect 4470 53 4544 57
<< metal3 >>
rect 260 253 387 513
rect 347 100 387 253
rect 4628 499 4654 500
rect 4628 490 4644 499
rect 4653 490 4654 499
rect 4628 489 4654 490
rect 347 99 488 100
rect 347 65 413 99
rect 487 65 488 99
rect 347 64 488 65
rect 4628 59 4638 489
rect 4468 57 4638 59
rect 4468 53 4470 57
rect 4544 53 4638 57
rect 4468 51 4638 53
use bondingpad  bondingpad_1
timestamp 1259953556
transform 1 0 0 0 -1 513
box 0 0 260 260
use bondingpad  bondingpad_0
timestamp 1259953556
transform 1 0 4740 0 -1 513
box 0 0 260 260
<< labels >>
rlabel m2contact 4307 0 4307 0 8 Gnd
rlabel m2contact 4441 0 4441 0 8 CVdd
rlabel m2contact 4412 0 4412 0 8 Bias
rlabel m2contact 4379 0 4379 0 8 Bias
rlabel m2contact 4351 0 4351 0 8 CVdd
rlabel m2contact 3833 0 3833 0 8 Gnd
rlabel m2contact 4011 0 4011 0 8 Gnd
rlabel m2contact 3967 0 3967 0 8 CVdd
rlabel m2contact 3938 0 3938 0 8 Bias
rlabel m2contact 3905 0 3905 0 8 Bias
rlabel m2contact 3877 0 3877 0 8 CVdd
rlabel m2contact 3359 0 3359 0 8 Gnd
rlabel m2contact 3537 0 3537 0 8 Gnd
rlabel m2contact 3493 0 3493 0 8 CVdd
rlabel m2contact 3464 0 3464 0 8 Bias
rlabel m2contact 3431 0 3431 0 8 Bias
rlabel m2contact 3403 0 3403 0 8 CVdd
rlabel m2contact 2885 0 2885 0 8 Gnd
rlabel m2contact 3063 0 3063 0 8 Gnd
rlabel m2contact 3019 0 3019 0 8 CVdd
rlabel m2contact 2990 0 2990 0 8 Bias
rlabel m2contact 2957 0 2957 0 8 Bias
rlabel m2contact 2929 0 2929 0 8 CVdd
rlabel m2contact 2411 0 2411 0 8 Gnd
rlabel m2contact 2589 0 2589 0 8 Gnd
rlabel m2contact 2545 0 2545 0 8 CVdd
rlabel m2contact 2516 0 2516 0 8 Bias
rlabel m2contact 2483 0 2483 0 8 Bias
rlabel m2contact 2455 0 2455 0 8 CVdd
rlabel m2contact 1937 0 1937 0 8 Gnd
rlabel m2contact 2115 0 2115 0 8 Gnd
rlabel m2contact 2071 0 2071 0 8 CVdd
rlabel m2contact 2042 0 2042 0 8 Bias
rlabel m2contact 2009 0 2009 0 8 Bias
rlabel m2contact 1981 0 1981 0 8 CVdd
rlabel m2contact 1463 0 1463 0 8 Gnd
rlabel m2contact 1641 0 1641 0 8 Gnd
rlabel m2contact 1597 0 1597 0 8 CVdd
rlabel m2contact 1568 0 1568 0 8 Bias
rlabel m2contact 1535 0 1535 0 8 Bias
rlabel m2contact 1507 0 1507 0 8 CVdd
rlabel m2contact 989 0 989 0 8 Gnd
rlabel m2contact 1167 0 1167 0 8 Gnd
rlabel m2contact 1123 0 1123 0 8 CVdd
rlabel m2contact 1094 0 1094 0 8 Bias
rlabel m2contact 1061 0 1061 0 8 Bias
rlabel m2contact 1033 0 1033 0 8 CVdd
rlabel m2contact 693 0 693 0 8 Gnd
rlabel m2contact 649 0 649 0 8 CVdd
rlabel m2contact 620 0 620 0 8 Bias
rlabel m2contact 587 0 587 0 8 Bias
rlabel m2contact 559 0 559 0 8 CVdd
<< end >>
