magic
tech scmos
timestamp 1418847243
<< nwell >>
rect 0 262 99 279
rect 0 168 99 210
rect -5 134 108 168
rect -26 83 -10 107
rect -10 51 108 60
rect -26 27 108 51
rect -5 16 108 27
<< pwell >>
rect 0 210 99 262
rect -5 89 108 134
rect -10 83 108 89
rect -26 70 108 83
rect -26 51 -10 70
rect -5 -21 108 10
<< psubstratepcontact >>
rect 3 242 7 246
rect 23 242 27 246
rect 47 242 51 246
rect 71 242 75 246
rect -2 117 2 121
rect 25 117 29 121
rect 52 117 56 121
rect 79 117 83 121
rect -2 -7 2 -3
rect 25 -7 29 -3
rect 52 -7 56 -3
rect 79 -7 83 -3
<< nsubstratencontact >>
rect 23 268 27 272
rect 47 268 51 272
rect 71 268 75 272
rect -2 150 2 154
rect 25 150 29 154
rect 52 150 56 154
rect 79 150 83 154
rect -2 26 2 30
rect 25 26 29 30
rect 52 26 56 30
rect 79 26 83 30
<< polysilicon >>
rect -12 231 2 233
rect -10 155 0 157
rect -10 89 -8 155
rect -10 81 0 89
rect -10 77 -8 81
rect -10 75 -3 77
rect -14 62 -11 64
rect -5 49 -3 75
rect -10 47 0 49
rect -10 -8 -8 47
rect -10 -10 0 -8
<< polycontact >>
rect -16 229 -12 233
rect -2 173 2 177
rect -4 93 0 97
rect -27 81 -23 85
rect -13 58 -9 62
rect -27 49 -23 53
<< metal1 >>
rect 3 275 83 279
rect 3 272 7 275
rect 23 272 27 275
rect 31 272 35 275
rect 47 272 51 275
rect 55 272 59 275
rect 71 272 75 275
rect 79 272 83 275
rect -3 268 8 272
rect 3 246 7 256
rect 0 237 3 245
rect 23 252 31 256
rect 47 252 55 256
rect 71 252 79 256
rect 23 246 27 252
rect 47 246 51 252
rect 71 246 75 252
rect 24 237 27 242
rect 48 237 51 242
rect 72 237 75 242
rect 0 233 2 237
rect -7 189 2 193
rect -16 173 -2 177
rect -7 158 1 161
rect -7 157 2 158
rect -2 154 2 157
rect 25 154 29 157
rect 52 154 56 159
rect 79 154 83 160
rect -14 97 -11 101
rect -4 85 0 93
rect -14 81 0 85
rect -14 65 -4 69
rect -9 58 0 61
rect -3 53 3 54
rect -14 51 3 53
rect -14 49 0 51
rect -14 33 -11 37
rect -7 30 3 34
rect -2 -10 2 -7
rect 25 -10 29 -7
rect 52 -10 56 -7
rect 79 -10 83 -7
<< m2contact >>
rect -7 268 -3 272
rect -4 233 0 237
rect -20 229 -16 233
rect -11 189 -7 193
rect -20 173 -16 177
rect 6 165 10 169
rect 17 165 21 169
rect 30 165 34 169
rect 41 165 45 169
rect 54 165 58 169
rect 65 165 69 169
rect 78 165 82 169
rect 89 165 93 169
rect -11 157 -7 161
rect -4 113 0 117
rect -11 97 -7 101
rect -20 81 -16 85
rect -4 65 0 69
rect -11 30 -7 37
rect -4 -14 0 -10
<< metal2 >>
rect -20 177 -17 229
rect -11 193 -7 272
rect -20 85 -17 173
rect -11 161 -7 189
rect -11 101 -7 157
rect -11 37 -7 97
rect -4 117 0 233
rect 6 136 10 165
rect 17 136 21 165
rect 30 132 34 165
rect 41 132 45 165
rect 69 165 75 169
rect 54 136 58 165
rect 71 136 75 165
rect 93 165 102 169
rect 78 136 82 165
rect 98 136 102 165
rect 54 132 62 136
rect 71 132 73 136
rect 78 132 87 136
rect -4 69 0 113
rect -4 -10 0 65
use dflipflopsimple  dflipflopsimple_0
array 0 3 24 0 0 76
timestamp 1418846892
transform -1 0 88 0 -1 88
box -10 -186 14 -81
use inverter  inverter_1
timestamp 1417997274
transform 1 0 -20 0 1 70
box -3 -5 6 31
use invinverter  invinverter_0
timestamp 1418010646
transform 1 0 -19 0 1 38
box -4 -5 5 31
use dflipflop  dflipflop_0
array 0 3 27 0 0 161
timestamp 1418018074
transform 1 0 11 0 1 135
box -11 -150 16 27
<< labels >>
rlabel metal2 -4 0 0 4 1 Gnd
rlabel m2contact -11 189 -7 193 1 Vdd
<< end >>
