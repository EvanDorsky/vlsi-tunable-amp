magic
tech scmos
timestamp 1418878488
<< nwell >>
rect -618 -4 0 117
rect 58 0 62 3
rect 43 -4 86 0
rect 141 0 150 7
rect 172 0 790 120
rect 129 -4 790 0
rect -618 -136 2 -4
rect 58 -5 62 -4
rect 141 -9 145 -4
rect 153 -5 157 -4
rect 172 -136 790 -4
<< pwell >>
rect 0 -4 43 3
rect 86 -4 129 3
rect -618 -378 2 -136
rect 5 -378 9 -268
rect 165 -378 169 -269
rect 172 -378 790 -136
rect -618 -393 790 -378
rect -4 -394 790 -393
<< electrodecontact >>
rect -626 -130 -622 22
rect 793 -124 797 26
<< electrodecap >>
rect -776 -132 -620 24
rect 791 -128 947 28
<< ntransistor >>
rect -606 -387 -600 -147
rect -594 -387 -588 -147
rect -582 -387 -576 -147
rect -570 -387 -564 -147
rect -558 -387 -552 -147
rect -546 -387 -540 -147
rect -534 -387 -528 -147
rect -522 -387 -516 -147
rect -510 -387 -504 -147
rect -498 -387 -492 -147
rect -486 -387 -480 -147
rect -474 -387 -468 -147
rect -462 -387 -456 -147
rect -450 -387 -444 -147
rect -438 -387 -432 -147
rect -426 -387 -420 -147
rect -414 -387 -408 -147
rect -402 -387 -396 -147
rect -390 -387 -384 -147
rect -378 -387 -372 -147
rect -366 -387 -360 -147
rect -354 -387 -348 -147
rect -342 -387 -336 -147
rect -330 -387 -324 -147
rect -318 -387 -312 -147
rect -306 -387 -300 -147
rect -294 -387 -288 -147
rect -282 -387 -276 -147
rect -270 -387 -264 -147
rect -258 -387 -252 -147
rect -246 -387 -240 -147
rect -234 -387 -228 -147
rect -222 -387 -216 -147
rect -210 -387 -204 -147
rect -198 -387 -192 -147
rect -186 -387 -180 -147
rect -174 -387 -168 -147
rect -162 -387 -156 -147
rect -150 -387 -144 -147
rect -138 -387 -132 -147
rect -126 -387 -120 -147
rect -114 -387 -108 -147
rect -102 -387 -96 -147
rect -90 -387 -84 -147
rect -78 -387 -72 -147
rect -66 -387 -60 -147
rect -54 -387 -48 -147
rect -42 -387 -36 -147
rect -30 -387 -24 -147
rect -18 -387 -12 -147
rect 184 -387 190 -147
rect 196 -387 202 -147
rect 208 -387 214 -147
rect 220 -387 226 -147
rect 232 -387 238 -147
rect 244 -387 250 -147
rect 256 -387 262 -147
rect 268 -387 274 -147
rect 280 -387 286 -147
rect 292 -387 298 -147
rect 304 -387 310 -147
rect 316 -387 322 -147
rect 328 -387 334 -147
rect 340 -387 346 -147
rect 352 -387 358 -147
rect 364 -387 370 -147
rect 376 -387 382 -147
rect 388 -387 394 -147
rect 400 -387 406 -147
rect 412 -387 418 -147
rect 424 -387 430 -147
rect 436 -387 442 -147
rect 448 -387 454 -147
rect 460 -387 466 -147
rect 472 -387 478 -147
rect 484 -387 490 -147
rect 496 -387 502 -147
rect 508 -387 514 -147
rect 520 -387 526 -147
rect 532 -387 538 -147
rect 544 -387 550 -147
rect 556 -387 562 -147
rect 568 -387 574 -147
rect 580 -387 586 -147
rect 592 -387 598 -147
rect 604 -387 610 -147
rect 616 -387 622 -147
rect 628 -387 634 -147
rect 640 -387 646 -147
rect 652 -387 658 -147
rect 664 -387 670 -147
rect 676 -387 682 -147
rect 688 -387 694 -147
rect 700 -387 706 -147
rect 712 -387 718 -147
rect 724 -387 730 -147
rect 736 -387 742 -147
rect 748 -387 754 -147
rect 760 -387 766 -147
rect 772 -387 778 -147
<< ptransistor >>
rect -606 -129 -600 111
rect -594 -129 -588 111
rect -582 -129 -576 111
rect -570 -129 -564 111
rect -558 -129 -552 111
rect -546 -129 -540 111
rect -534 -129 -528 111
rect -522 -129 -516 111
rect -510 -129 -504 111
rect -498 -129 -492 111
rect -486 -129 -480 111
rect -474 -129 -468 111
rect -462 -129 -456 111
rect -450 -129 -444 111
rect -438 -129 -432 111
rect -426 -129 -420 111
rect -414 -129 -408 111
rect -402 -129 -396 111
rect -390 -129 -384 111
rect -378 -129 -372 111
rect -366 -129 -360 111
rect -354 -129 -348 111
rect -342 -129 -336 111
rect -330 -129 -324 111
rect -318 -129 -312 111
rect -306 -129 -300 111
rect -294 -129 -288 111
rect -282 -129 -276 111
rect -270 -129 -264 111
rect -258 -129 -252 111
rect -246 -129 -240 111
rect -234 -129 -228 111
rect -222 -129 -216 111
rect -210 -129 -204 111
rect -198 -129 -192 111
rect -186 -129 -180 111
rect -174 -129 -168 111
rect -162 -129 -156 111
rect -150 -129 -144 111
rect -138 -129 -132 111
rect -126 -129 -120 111
rect -114 -129 -108 111
rect -102 -129 -96 111
rect -90 -129 -84 111
rect -78 -129 -72 111
rect -66 -129 -60 111
rect -54 -129 -48 111
rect -42 -129 -36 111
rect -30 -129 -24 111
rect -18 -129 -12 111
rect 184 -126 190 114
rect 196 -126 202 114
rect 208 -126 214 114
rect 220 -126 226 114
rect 232 -126 238 114
rect 244 -126 250 114
rect 256 -126 262 114
rect 268 -126 274 114
rect 280 -126 286 114
rect 292 -126 298 114
rect 304 -126 310 114
rect 316 -126 322 114
rect 328 -126 334 114
rect 340 -126 346 114
rect 352 -126 358 114
rect 364 -126 370 114
rect 376 -126 382 114
rect 388 -126 394 114
rect 400 -126 406 114
rect 412 -126 418 114
rect 424 -126 430 114
rect 436 -126 442 114
rect 448 -126 454 114
rect 460 -126 466 114
rect 472 -126 478 114
rect 484 -126 490 114
rect 496 -126 502 114
rect 508 -126 514 114
rect 520 -126 526 114
rect 532 -126 538 114
rect 544 -126 550 114
rect 556 -126 562 114
rect 568 -126 574 114
rect 580 -126 586 114
rect 592 -126 598 114
rect 604 -126 610 114
rect 616 -126 622 114
rect 628 -126 634 114
rect 640 -126 646 114
rect 652 -126 658 114
rect 664 -126 670 114
rect 676 -126 682 114
rect 688 -126 694 114
rect 700 -126 706 114
rect 712 -126 718 114
rect 724 -126 730 114
rect 736 -126 742 114
rect 748 -126 754 114
rect 760 -126 766 114
rect 772 -126 778 114
<< ndiffusion >>
rect -612 -387 -611 -147
rect -607 -387 -606 -147
rect -600 -387 -599 -147
rect -595 -387 -594 -147
rect -588 -387 -587 -147
rect -583 -387 -582 -147
rect -576 -387 -575 -147
rect -571 -387 -570 -147
rect -564 -387 -563 -147
rect -559 -387 -558 -147
rect -552 -387 -551 -147
rect -547 -387 -546 -147
rect -540 -387 -539 -147
rect -535 -387 -534 -147
rect -528 -387 -527 -147
rect -523 -387 -522 -147
rect -516 -387 -515 -147
rect -511 -387 -510 -147
rect -504 -387 -503 -147
rect -499 -387 -498 -147
rect -492 -387 -491 -147
rect -487 -387 -486 -147
rect -480 -387 -479 -147
rect -475 -387 -474 -147
rect -468 -387 -467 -147
rect -463 -387 -462 -147
rect -456 -387 -455 -147
rect -451 -387 -450 -147
rect -444 -387 -443 -147
rect -439 -387 -438 -147
rect -432 -387 -431 -147
rect -427 -387 -426 -147
rect -420 -387 -419 -147
rect -415 -387 -414 -147
rect -408 -387 -407 -147
rect -403 -387 -402 -147
rect -396 -387 -395 -147
rect -391 -387 -390 -147
rect -384 -387 -383 -147
rect -379 -387 -378 -147
rect -372 -387 -371 -147
rect -367 -387 -366 -147
rect -360 -387 -359 -147
rect -355 -387 -354 -147
rect -348 -387 -347 -147
rect -343 -387 -342 -147
rect -336 -387 -335 -147
rect -331 -387 -330 -147
rect -324 -387 -323 -147
rect -319 -387 -318 -147
rect -312 -387 -311 -147
rect -307 -387 -306 -147
rect -300 -387 -299 -147
rect -295 -387 -294 -147
rect -288 -387 -287 -147
rect -283 -387 -282 -147
rect -276 -387 -275 -147
rect -271 -387 -270 -147
rect -264 -387 -263 -147
rect -259 -387 -258 -147
rect -252 -387 -251 -147
rect -247 -387 -246 -147
rect -240 -387 -239 -147
rect -235 -387 -234 -147
rect -228 -387 -227 -147
rect -223 -387 -222 -147
rect -216 -387 -215 -147
rect -211 -387 -210 -147
rect -204 -387 -203 -147
rect -199 -387 -198 -147
rect -192 -387 -191 -147
rect -187 -387 -186 -147
rect -180 -387 -179 -147
rect -175 -387 -174 -147
rect -168 -387 -167 -147
rect -163 -387 -162 -147
rect -156 -387 -155 -147
rect -151 -387 -150 -147
rect -144 -387 -143 -147
rect -139 -387 -138 -147
rect -132 -387 -131 -147
rect -127 -387 -126 -147
rect -120 -387 -119 -147
rect -115 -387 -114 -147
rect -108 -387 -107 -147
rect -103 -387 -102 -147
rect -96 -387 -95 -147
rect -91 -387 -90 -147
rect -84 -387 -83 -147
rect -79 -387 -78 -147
rect -72 -387 -71 -147
rect -67 -387 -66 -147
rect -60 -387 -59 -147
rect -55 -387 -54 -147
rect -48 -387 -47 -147
rect -43 -387 -42 -147
rect -36 -387 -35 -147
rect -31 -387 -30 -147
rect -24 -387 -23 -147
rect -19 -387 -18 -147
rect -12 -387 -11 -147
rect -7 -387 -6 -147
rect 178 -387 179 -147
rect 183 -387 184 -147
rect 190 -387 191 -147
rect 195 -387 196 -147
rect 202 -387 203 -147
rect 207 -387 208 -147
rect 214 -387 215 -147
rect 219 -387 220 -147
rect 226 -387 227 -147
rect 231 -387 232 -147
rect 238 -387 239 -147
rect 243 -387 244 -147
rect 250 -387 251 -147
rect 255 -387 256 -147
rect 262 -387 263 -147
rect 267 -387 268 -147
rect 274 -387 275 -147
rect 279 -387 280 -147
rect 286 -387 287 -147
rect 291 -387 292 -147
rect 298 -387 299 -147
rect 303 -387 304 -147
rect 310 -387 311 -147
rect 315 -387 316 -147
rect 322 -387 323 -147
rect 327 -387 328 -147
rect 334 -387 335 -147
rect 339 -387 340 -147
rect 346 -387 347 -147
rect 351 -387 352 -147
rect 358 -387 359 -147
rect 363 -387 364 -147
rect 370 -387 371 -147
rect 375 -387 376 -147
rect 382 -387 383 -147
rect 387 -387 388 -147
rect 394 -387 395 -147
rect 399 -387 400 -147
rect 406 -387 407 -147
rect 411 -387 412 -147
rect 418 -387 419 -147
rect 423 -387 424 -147
rect 430 -387 431 -147
rect 435 -387 436 -147
rect 442 -387 443 -147
rect 447 -387 448 -147
rect 454 -387 455 -147
rect 459 -387 460 -147
rect 466 -387 467 -147
rect 471 -387 472 -147
rect 478 -387 479 -147
rect 483 -387 484 -147
rect 490 -387 491 -147
rect 495 -387 496 -147
rect 502 -387 503 -147
rect 507 -387 508 -147
rect 514 -387 515 -147
rect 519 -387 520 -147
rect 526 -387 527 -147
rect 531 -387 532 -147
rect 538 -387 539 -147
rect 543 -387 544 -147
rect 550 -387 551 -147
rect 555 -387 556 -147
rect 562 -387 563 -147
rect 567 -387 568 -147
rect 574 -387 575 -147
rect 579 -387 580 -147
rect 586 -387 587 -147
rect 591 -387 592 -147
rect 598 -387 599 -147
rect 603 -387 604 -147
rect 610 -387 611 -147
rect 615 -387 616 -147
rect 622 -387 623 -147
rect 627 -387 628 -147
rect 634 -387 635 -147
rect 639 -387 640 -147
rect 646 -387 647 -147
rect 651 -387 652 -147
rect 658 -387 659 -147
rect 663 -387 664 -147
rect 670 -387 671 -147
rect 675 -387 676 -147
rect 682 -387 683 -147
rect 687 -387 688 -147
rect 694 -387 695 -147
rect 699 -387 700 -147
rect 706 -387 707 -147
rect 711 -387 712 -147
rect 718 -387 719 -147
rect 723 -387 724 -147
rect 730 -387 731 -147
rect 735 -387 736 -147
rect 742 -387 743 -147
rect 747 -387 748 -147
rect 754 -387 755 -147
rect 759 -387 760 -147
rect 766 -387 767 -147
rect 771 -387 772 -147
rect 778 -387 779 -147
rect 783 -387 784 -147
<< pdiffusion >>
rect -612 -129 -611 111
rect -607 -129 -606 111
rect -600 -129 -599 111
rect -595 -129 -594 111
rect -588 -129 -587 111
rect -583 -129 -582 111
rect -576 -129 -575 111
rect -571 -129 -570 111
rect -564 -129 -563 111
rect -559 -129 -558 111
rect -552 -129 -551 111
rect -547 -129 -546 111
rect -540 -129 -539 111
rect -535 -129 -534 111
rect -528 -129 -527 111
rect -523 -129 -522 111
rect -516 -129 -515 111
rect -511 -129 -510 111
rect -504 -129 -503 111
rect -499 -129 -498 111
rect -492 -129 -491 111
rect -487 -129 -486 111
rect -480 -129 -479 111
rect -475 -129 -474 111
rect -468 -129 -467 111
rect -463 -129 -462 111
rect -456 -129 -455 111
rect -451 -129 -450 111
rect -444 -129 -443 111
rect -439 -129 -438 111
rect -432 -129 -431 111
rect -427 -129 -426 111
rect -420 -129 -419 111
rect -415 -129 -414 111
rect -408 -129 -407 111
rect -403 -129 -402 111
rect -396 -129 -395 111
rect -391 -129 -390 111
rect -384 -129 -383 111
rect -379 -129 -378 111
rect -372 -129 -371 111
rect -367 -129 -366 111
rect -360 -129 -359 111
rect -355 -129 -354 111
rect -348 -129 -347 111
rect -343 -129 -342 111
rect -336 -129 -335 111
rect -331 -129 -330 111
rect -324 -129 -323 111
rect -319 -129 -318 111
rect -312 -129 -311 111
rect -307 -129 -306 111
rect -300 -129 -299 111
rect -295 -129 -294 111
rect -288 -129 -287 111
rect -283 -129 -282 111
rect -276 -129 -275 111
rect -271 -129 -270 111
rect -264 -129 -263 111
rect -259 -129 -258 111
rect -252 -129 -251 111
rect -247 -129 -246 111
rect -240 -129 -239 111
rect -235 -129 -234 111
rect -228 -129 -227 111
rect -223 -129 -222 111
rect -216 -129 -215 111
rect -211 -129 -210 111
rect -204 -129 -203 111
rect -199 -129 -198 111
rect -192 -129 -191 111
rect -187 -129 -186 111
rect -180 -129 -179 111
rect -175 -129 -174 111
rect -168 -129 -167 111
rect -163 -129 -162 111
rect -156 -129 -155 111
rect -151 -129 -150 111
rect -144 -129 -143 111
rect -139 -129 -138 111
rect -132 -129 -131 111
rect -127 -129 -126 111
rect -120 -129 -119 111
rect -115 -129 -114 111
rect -108 -129 -107 111
rect -103 -129 -102 111
rect -96 -129 -95 111
rect -91 -129 -90 111
rect -84 -129 -83 111
rect -79 -129 -78 111
rect -72 -129 -71 111
rect -67 -129 -66 111
rect -60 -129 -59 111
rect -55 -129 -54 111
rect -48 -129 -47 111
rect -43 -129 -42 111
rect -36 -129 -35 111
rect -31 -129 -30 111
rect -24 -129 -23 111
rect -19 -129 -18 111
rect -12 -129 -11 111
rect -7 -129 -6 111
rect 178 -126 179 114
rect 183 -126 184 114
rect 190 -126 191 114
rect 195 -126 196 114
rect 202 -126 203 114
rect 207 -126 208 114
rect 214 -126 215 114
rect 219 -126 220 114
rect 226 -126 227 114
rect 231 -126 232 114
rect 238 -126 239 114
rect 243 -126 244 114
rect 250 -126 251 114
rect 255 -126 256 114
rect 262 -126 263 114
rect 267 -126 268 114
rect 274 -126 275 114
rect 279 -126 280 114
rect 286 -126 287 114
rect 291 -126 292 114
rect 298 -126 299 114
rect 303 -126 304 114
rect 310 -126 311 114
rect 315 -126 316 114
rect 322 -126 323 114
rect 327 -126 328 114
rect 334 -126 335 114
rect 339 -126 340 114
rect 346 -126 347 114
rect 351 -126 352 114
rect 358 -126 359 114
rect 363 -126 364 114
rect 370 -126 371 114
rect 375 -126 376 114
rect 382 -126 383 114
rect 387 -126 388 114
rect 394 -126 395 114
rect 399 -126 400 114
rect 406 -126 407 114
rect 411 -126 412 114
rect 418 -126 419 114
rect 423 -126 424 114
rect 430 -126 431 114
rect 435 -126 436 114
rect 442 -126 443 114
rect 447 -126 448 114
rect 454 -126 455 114
rect 459 -126 460 114
rect 466 -126 467 114
rect 471 -126 472 114
rect 478 -126 479 114
rect 483 -126 484 114
rect 490 -126 491 114
rect 495 -126 496 114
rect 502 -126 503 114
rect 507 -126 508 114
rect 514 -126 515 114
rect 519 -126 520 114
rect 526 -126 527 114
rect 531 -126 532 114
rect 538 -126 539 114
rect 543 -126 544 114
rect 550 -126 551 114
rect 555 -126 556 114
rect 562 -126 563 114
rect 567 -126 568 114
rect 574 -126 575 114
rect 579 -126 580 114
rect 586 -126 587 114
rect 591 -126 592 114
rect 598 -126 599 114
rect 603 -126 604 114
rect 610 -126 611 114
rect 615 -126 616 114
rect 622 -126 623 114
rect 627 -126 628 114
rect 634 -126 635 114
rect 639 -126 640 114
rect 646 -126 647 114
rect 651 -126 652 114
rect 658 -126 659 114
rect 663 -126 664 114
rect 670 -126 671 114
rect 675 -126 676 114
rect 682 -126 683 114
rect 687 -126 688 114
rect 694 -126 695 114
rect 699 -126 700 114
rect 706 -126 707 114
rect 711 -126 712 114
rect 718 -126 719 114
rect 723 -126 724 114
rect 730 -126 731 114
rect 735 -126 736 114
rect 742 -126 743 114
rect 747 -126 748 114
rect 754 -126 755 114
rect 759 -126 760 114
rect 766 -126 767 114
rect 771 -126 772 114
rect 778 -126 779 114
rect 783 -126 784 114
<< ndcontact >>
rect -611 -387 -607 -147
rect -599 -387 -595 -147
rect -587 -387 -583 -147
rect -575 -387 -571 -147
rect -563 -387 -559 -147
rect -551 -387 -547 -147
rect -539 -387 -535 -147
rect -527 -387 -523 -147
rect -515 -387 -511 -147
rect -503 -387 -499 -147
rect -491 -387 -487 -147
rect -479 -387 -475 -147
rect -467 -387 -463 -147
rect -455 -387 -451 -147
rect -443 -387 -439 -147
rect -431 -387 -427 -147
rect -419 -387 -415 -147
rect -407 -387 -403 -147
rect -395 -387 -391 -147
rect -383 -387 -379 -147
rect -371 -387 -367 -147
rect -359 -387 -355 -147
rect -347 -387 -343 -147
rect -335 -387 -331 -147
rect -323 -387 -319 -147
rect -311 -387 -307 -147
rect -299 -387 -295 -147
rect -287 -387 -283 -147
rect -275 -387 -271 -147
rect -263 -387 -259 -147
rect -251 -387 -247 -147
rect -239 -387 -235 -147
rect -227 -387 -223 -147
rect -215 -387 -211 -147
rect -203 -387 -199 -147
rect -191 -387 -187 -147
rect -179 -387 -175 -147
rect -167 -387 -163 -147
rect -155 -387 -151 -147
rect -143 -387 -139 -147
rect -131 -387 -127 -147
rect -119 -387 -115 -147
rect -107 -387 -103 -147
rect -95 -387 -91 -147
rect -83 -387 -79 -147
rect -71 -387 -67 -147
rect -59 -387 -55 -147
rect -47 -387 -43 -147
rect -35 -387 -31 -147
rect -23 -387 -19 -147
rect -11 -387 -7 -147
rect 179 -387 183 -147
rect 191 -387 195 -147
rect 203 -387 207 -147
rect 215 -387 219 -147
rect 227 -387 231 -147
rect 239 -387 243 -147
rect 251 -387 255 -147
rect 263 -387 267 -147
rect 275 -387 279 -147
rect 287 -387 291 -147
rect 299 -387 303 -147
rect 311 -387 315 -147
rect 323 -387 327 -147
rect 335 -387 339 -147
rect 347 -387 351 -147
rect 359 -387 363 -147
rect 371 -387 375 -147
rect 383 -387 387 -147
rect 395 -387 399 -147
rect 407 -387 411 -147
rect 419 -387 423 -147
rect 431 -387 435 -147
rect 443 -387 447 -147
rect 455 -387 459 -147
rect 467 -387 471 -147
rect 479 -387 483 -147
rect 491 -387 495 -147
rect 503 -387 507 -147
rect 515 -387 519 -147
rect 527 -387 531 -147
rect 539 -387 543 -147
rect 551 -387 555 -147
rect 563 -387 567 -147
rect 575 -387 579 -147
rect 587 -387 591 -147
rect 599 -387 603 -147
rect 611 -387 615 -147
rect 623 -387 627 -147
rect 635 -387 639 -147
rect 647 -387 651 -147
rect 659 -387 663 -147
rect 671 -387 675 -147
rect 683 -387 687 -147
rect 695 -387 699 -147
rect 707 -387 711 -147
rect 719 -387 723 -147
rect 731 -387 735 -147
rect 743 -387 747 -147
rect 755 -387 759 -147
rect 767 -387 771 -147
rect 779 -387 783 -147
<< pdcontact >>
rect -611 -129 -607 111
rect -599 -129 -595 111
rect -587 -129 -583 111
rect -575 -129 -571 111
rect -563 -129 -559 111
rect -551 -129 -547 111
rect -539 -129 -535 111
rect -527 -129 -523 111
rect -515 -129 -511 111
rect -503 -129 -499 111
rect -491 -129 -487 111
rect -479 -129 -475 111
rect -467 -129 -463 111
rect -455 -129 -451 111
rect -443 -129 -439 111
rect -431 -129 -427 111
rect -419 -129 -415 111
rect -407 -129 -403 111
rect -395 -129 -391 111
rect -383 -129 -379 111
rect -371 -129 -367 111
rect -359 -129 -355 111
rect -347 -129 -343 111
rect -335 -129 -331 111
rect -323 -129 -319 111
rect -311 -129 -307 111
rect -299 -129 -295 111
rect -287 -129 -283 111
rect -275 -129 -271 111
rect -263 -129 -259 111
rect -251 -129 -247 111
rect -239 -129 -235 111
rect -227 -129 -223 111
rect -215 -129 -211 111
rect -203 -129 -199 111
rect -191 -129 -187 111
rect -179 -129 -175 111
rect -167 -129 -163 111
rect -155 -129 -151 111
rect -143 -129 -139 111
rect -131 -129 -127 111
rect -119 -129 -115 111
rect -107 -129 -103 111
rect -95 -129 -91 111
rect -83 -129 -79 111
rect -71 -129 -67 111
rect -59 -129 -55 111
rect -47 -129 -43 111
rect -35 -129 -31 111
rect -23 -129 -19 111
rect -11 -129 -7 111
rect 11 -14 15 -10
rect 103 -14 107 -10
rect 179 -126 183 114
rect 191 -126 195 114
rect 203 -126 207 114
rect 215 -126 219 114
rect 227 -126 231 114
rect 239 -126 243 114
rect 251 -126 255 114
rect 263 -126 267 114
rect 275 -126 279 114
rect 287 -126 291 114
rect 299 -126 303 114
rect 311 -126 315 114
rect 323 -126 327 114
rect 335 -126 339 114
rect 347 -126 351 114
rect 359 -126 363 114
rect 371 -126 375 114
rect 383 -126 387 114
rect 395 -126 399 114
rect 407 -126 411 114
rect 419 -126 423 114
rect 431 -126 435 114
rect 443 -126 447 114
rect 455 -126 459 114
rect 467 -126 471 114
rect 479 -126 483 114
rect 491 -126 495 114
rect 503 -126 507 114
rect 515 -126 519 114
rect 527 -126 531 114
rect 539 -126 543 114
rect 551 -126 555 114
rect 563 -126 567 114
rect 575 -126 579 114
rect 587 -126 591 114
rect 599 -126 603 114
rect 611 -126 615 114
rect 623 -126 627 114
rect 635 -126 639 114
rect 647 -126 651 114
rect 659 -126 663 114
rect 671 -126 675 114
rect 683 -126 687 114
rect 695 -126 699 114
rect 707 -126 711 114
rect 719 -126 723 114
rect 731 -126 735 114
rect 743 -126 747 114
rect 755 -126 759 114
rect 767 -126 771 114
rect 779 -126 783 114
<< psubstratepcontact >>
rect 5 -383 9 -268
rect 165 -383 169 -269
<< polysilicon >>
rect 185 119 189 124
rect -606 114 -15 116
rect 184 115 778 119
rect 184 114 190 115
rect 196 114 202 115
rect 208 114 214 115
rect 220 114 226 115
rect 232 114 238 115
rect 244 114 250 115
rect 256 114 262 115
rect 268 114 274 115
rect 280 114 286 115
rect 292 114 298 115
rect 304 114 310 115
rect 316 114 322 115
rect 328 114 334 115
rect 340 114 346 115
rect 352 114 358 115
rect 364 114 370 115
rect 376 114 382 115
rect 388 114 394 115
rect 400 114 406 115
rect 412 114 418 115
rect 424 114 430 115
rect 436 114 442 115
rect 448 114 454 115
rect 460 114 466 115
rect 472 114 478 115
rect 484 114 490 115
rect 496 114 502 115
rect 508 114 514 115
rect 520 114 526 115
rect 532 114 538 115
rect 544 114 550 115
rect 556 114 562 115
rect 568 114 574 115
rect 580 114 586 115
rect 592 114 598 115
rect 604 114 610 115
rect 616 114 622 115
rect 628 114 634 115
rect 640 114 646 115
rect 652 114 658 115
rect 664 114 670 115
rect 676 114 682 115
rect 688 114 694 115
rect 700 114 706 115
rect 712 114 718 115
rect 724 114 730 115
rect 736 114 742 115
rect 748 114 754 115
rect 760 114 766 115
rect 772 114 778 115
rect -606 112 -12 114
rect -606 111 -600 112
rect -594 111 -588 112
rect -582 111 -576 112
rect -570 111 -564 112
rect -558 111 -552 112
rect -546 111 -540 112
rect -534 111 -528 112
rect -522 111 -516 112
rect -510 111 -504 112
rect -498 111 -492 112
rect -486 111 -480 112
rect -474 111 -468 112
rect -462 111 -456 112
rect -450 111 -444 112
rect -438 111 -432 112
rect -426 111 -420 112
rect -414 111 -408 112
rect -402 111 -396 112
rect -390 111 -384 112
rect -378 111 -372 112
rect -366 111 -360 112
rect -354 111 -348 112
rect -342 111 -336 112
rect -330 111 -324 112
rect -318 111 -312 112
rect -306 111 -300 112
rect -294 111 -288 112
rect -282 111 -276 112
rect -270 111 -264 112
rect -258 111 -252 112
rect -246 111 -240 112
rect -234 111 -228 112
rect -222 111 -216 112
rect -210 111 -204 112
rect -198 111 -192 112
rect -186 111 -180 112
rect -174 111 -168 112
rect -162 111 -156 112
rect -150 111 -144 112
rect -138 111 -132 112
rect -126 111 -120 112
rect -114 111 -108 112
rect -102 111 -96 112
rect -90 111 -84 112
rect -78 111 -72 112
rect -66 111 -60 112
rect -54 111 -48 112
rect -42 111 -36 112
rect -30 111 -24 112
rect -18 111 -12 112
rect -781 -132 -615 29
rect 57 3 63 4
rect 109 3 115 4
rect 140 3 146 4
rect 184 -129 190 -126
rect 196 -129 202 -126
rect 208 -129 214 -126
rect 220 -129 226 -126
rect 232 -129 238 -126
rect 244 -129 250 -126
rect 256 -129 262 -126
rect 268 -129 274 -126
rect 280 -129 286 -126
rect 292 -129 298 -126
rect 304 -129 310 -126
rect 316 -129 322 -126
rect 328 -129 334 -126
rect 340 -129 346 -126
rect 352 -129 358 -126
rect 364 -129 370 -126
rect 376 -129 382 -126
rect 388 -129 394 -126
rect 400 -129 406 -126
rect 412 -129 418 -126
rect 424 -129 430 -126
rect 436 -129 442 -126
rect 448 -129 454 -126
rect 460 -129 466 -126
rect 472 -129 478 -126
rect 484 -129 490 -126
rect 496 -129 502 -126
rect 508 -129 514 -126
rect 520 -129 526 -126
rect 532 -129 538 -126
rect 544 -129 550 -126
rect 556 -129 562 -126
rect 568 -129 574 -126
rect 580 -129 586 -126
rect 592 -129 598 -126
rect 604 -129 610 -126
rect 616 -129 622 -126
rect 628 -129 634 -126
rect 640 -129 646 -126
rect 652 -129 658 -126
rect 664 -129 670 -126
rect 676 -129 682 -126
rect 688 -129 694 -126
rect 700 -129 706 -126
rect 712 -129 718 -126
rect 724 -129 730 -126
rect 736 -129 742 -126
rect 748 -129 754 -126
rect 760 -129 766 -126
rect 772 -129 778 -126
rect 786 -129 952 33
rect -606 -132 -600 -129
rect -594 -132 -588 -129
rect -582 -132 -576 -129
rect -570 -132 -564 -129
rect -558 -132 -552 -129
rect -546 -132 -540 -129
rect -534 -132 -528 -129
rect -522 -132 -516 -129
rect -510 -132 -504 -129
rect -498 -132 -492 -129
rect -486 -132 -480 -129
rect -474 -132 -468 -129
rect -462 -132 -456 -129
rect -450 -132 -444 -129
rect -438 -132 -432 -129
rect -426 -132 -420 -129
rect -414 -132 -408 -129
rect -402 -132 -396 -129
rect -390 -132 -384 -129
rect -378 -132 -372 -129
rect -366 -132 -360 -129
rect -354 -132 -348 -129
rect -342 -132 -336 -129
rect -330 -132 -324 -129
rect -318 -132 -312 -129
rect -306 -132 -300 -129
rect -294 -132 -288 -129
rect -282 -132 -276 -129
rect -270 -132 -264 -129
rect -258 -132 -252 -129
rect -246 -132 -240 -129
rect -234 -132 -228 -129
rect -222 -132 -216 -129
rect -210 -132 -204 -129
rect -198 -132 -192 -129
rect -186 -132 -180 -129
rect -174 -132 -168 -129
rect -162 -132 -156 -129
rect -150 -132 -144 -129
rect -138 -132 -132 -129
rect -126 -132 -120 -129
rect -114 -132 -108 -129
rect -102 -132 -96 -129
rect -90 -132 -84 -129
rect -78 -132 -72 -129
rect -66 -132 -60 -129
rect -54 -132 -48 -129
rect -42 -132 -36 -129
rect -30 -132 -24 -129
rect -18 -132 -12 -129
rect -781 -136 -12 -132
rect 179 -133 952 -129
rect -781 -137 -615 -136
rect -606 -144 -593 -142
rect -589 -144 -581 -142
rect -577 -144 -569 -142
rect -565 -144 -557 -142
rect -553 -144 -545 -142
rect -541 -144 -533 -142
rect -529 -144 -521 -142
rect -517 -144 -509 -142
rect -505 -144 -497 -142
rect -493 -144 -485 -142
rect -481 -144 -473 -142
rect -469 -144 -461 -142
rect -457 -144 -449 -142
rect -445 -144 -437 -142
rect -433 -144 -425 -142
rect -421 -144 -413 -142
rect -409 -144 -401 -142
rect -397 -144 -389 -142
rect -385 -144 -377 -142
rect -373 -144 -365 -142
rect -361 -144 -353 -142
rect -349 -144 -341 -142
rect -337 -144 -329 -142
rect -325 -144 -317 -142
rect -313 -144 -305 -142
rect -301 -144 -293 -142
rect -289 -144 -281 -142
rect -277 -144 -269 -142
rect -265 -144 -257 -142
rect -253 -144 -245 -142
rect -241 -144 -233 -142
rect -229 -144 -221 -142
rect -217 -144 -209 -142
rect -205 -144 -197 -142
rect -193 -144 -185 -142
rect -181 -144 -173 -142
rect -169 -144 -161 -142
rect -157 -144 -149 -142
rect -145 -144 -137 -142
rect -133 -144 -125 -142
rect -121 -144 -113 -142
rect -109 -144 -101 -142
rect -97 -144 -89 -142
rect -85 -144 -77 -142
rect -73 -144 -65 -142
rect -61 -144 -53 -142
rect -49 -144 -41 -142
rect -37 -144 -29 -142
rect -25 -144 -12 -142
rect -606 -146 -12 -144
rect -606 -147 -600 -146
rect -594 -147 -588 -146
rect -582 -147 -576 -146
rect -570 -147 -564 -146
rect -558 -147 -552 -146
rect -546 -147 -540 -146
rect -534 -147 -528 -146
rect -522 -147 -516 -146
rect -510 -147 -504 -146
rect -498 -147 -492 -146
rect -486 -147 -480 -146
rect -474 -147 -468 -146
rect -462 -147 -456 -146
rect -450 -147 -444 -146
rect -438 -147 -432 -146
rect -426 -147 -420 -146
rect -414 -147 -408 -146
rect -402 -147 -396 -146
rect -390 -147 -384 -146
rect -378 -147 -372 -146
rect -366 -147 -360 -146
rect -354 -147 -348 -146
rect -342 -147 -336 -146
rect -330 -147 -324 -146
rect -318 -147 -312 -146
rect -306 -147 -300 -146
rect -294 -147 -288 -146
rect -282 -147 -276 -146
rect -270 -147 -264 -146
rect -258 -147 -252 -146
rect -246 -147 -240 -146
rect -234 -147 -228 -146
rect -222 -147 -216 -146
rect -210 -147 -204 -146
rect -198 -147 -192 -146
rect -186 -147 -180 -146
rect -174 -147 -168 -146
rect -162 -147 -156 -146
rect -150 -147 -144 -146
rect -138 -147 -132 -146
rect -126 -147 -120 -146
rect -114 -147 -108 -146
rect -102 -147 -96 -146
rect -90 -147 -84 -146
rect -78 -147 -72 -146
rect -66 -147 -60 -146
rect -54 -147 -48 -146
rect -42 -147 -36 -146
rect -30 -147 -24 -146
rect -18 -147 -12 -146
rect 184 -146 778 -142
rect 184 -147 190 -146
rect 196 -147 202 -146
rect 208 -147 214 -146
rect 220 -147 226 -146
rect 232 -147 238 -146
rect 244 -147 250 -146
rect 256 -147 262 -146
rect 268 -147 274 -146
rect 280 -147 286 -146
rect 292 -147 298 -146
rect 304 -147 310 -146
rect 316 -147 322 -146
rect 328 -147 334 -146
rect 340 -147 346 -146
rect 352 -147 358 -146
rect 364 -147 370 -146
rect 376 -147 382 -146
rect 388 -147 394 -146
rect 400 -147 406 -146
rect 412 -147 418 -146
rect 424 -147 430 -146
rect 436 -147 442 -146
rect 448 -147 454 -146
rect 460 -147 466 -146
rect 472 -147 478 -146
rect 484 -147 490 -146
rect 496 -147 502 -146
rect 508 -147 514 -146
rect 520 -147 526 -146
rect 532 -147 538 -146
rect 544 -147 550 -146
rect 556 -147 562 -146
rect 568 -147 574 -146
rect 580 -147 586 -146
rect 592 -147 598 -146
rect 604 -147 610 -146
rect 616 -147 622 -146
rect 628 -147 634 -146
rect 640 -147 646 -146
rect 652 -147 658 -146
rect 664 -147 670 -146
rect 676 -147 682 -146
rect 688 -147 694 -146
rect 700 -147 706 -146
rect 712 -147 718 -146
rect 724 -147 730 -146
rect 736 -147 742 -146
rect 748 -147 754 -146
rect 760 -147 766 -146
rect 772 -147 778 -146
rect -606 -390 -600 -387
rect -594 -390 -588 -387
rect -582 -390 -576 -387
rect -570 -390 -564 -387
rect -558 -390 -552 -387
rect -546 -390 -540 -387
rect -534 -390 -528 -387
rect -522 -390 -516 -387
rect -510 -390 -504 -387
rect -498 -390 -492 -387
rect -486 -390 -480 -387
rect -474 -390 -468 -387
rect -462 -390 -456 -387
rect -450 -390 -444 -387
rect -438 -390 -432 -387
rect -426 -390 -420 -387
rect -414 -390 -408 -387
rect -402 -390 -396 -387
rect -390 -390 -384 -387
rect -378 -390 -372 -387
rect -366 -390 -360 -387
rect -354 -390 -348 -387
rect -342 -390 -336 -387
rect -330 -390 -324 -387
rect -318 -390 -312 -387
rect -306 -390 -300 -387
rect -294 -390 -288 -387
rect -282 -390 -276 -387
rect -270 -390 -264 -387
rect -258 -390 -252 -387
rect -246 -390 -240 -387
rect -234 -390 -228 -387
rect -222 -390 -216 -387
rect -210 -390 -204 -387
rect -198 -390 -192 -387
rect -186 -390 -180 -387
rect -174 -390 -168 -387
rect -162 -390 -156 -387
rect -150 -390 -144 -387
rect -138 -390 -132 -387
rect -126 -390 -120 -387
rect -114 -390 -108 -387
rect -102 -390 -96 -387
rect -90 -390 -84 -387
rect -78 -390 -72 -387
rect -66 -390 -60 -387
rect -54 -390 -48 -387
rect -42 -390 -36 -387
rect -30 -390 -24 -387
rect -18 -390 -12 -387
rect 184 -390 190 -387
rect 196 -390 202 -387
rect 208 -390 214 -387
rect 220 -390 226 -387
rect 232 -390 238 -387
rect 244 -390 250 -387
rect 256 -390 262 -387
rect 268 -390 274 -387
rect 280 -390 286 -387
rect 292 -390 298 -387
rect 304 -390 310 -387
rect 316 -390 322 -387
rect 328 -390 334 -387
rect 340 -390 346 -387
rect 352 -390 358 -387
rect 364 -390 370 -387
rect 376 -390 382 -387
rect 388 -390 394 -387
rect 400 -390 406 -387
rect 412 -390 418 -387
rect 424 -390 430 -387
rect 436 -390 442 -387
rect 448 -390 454 -387
rect 460 -390 466 -387
rect 472 -390 478 -387
rect 484 -390 490 -387
rect 496 -390 502 -387
rect 508 -390 514 -387
rect 520 -390 526 -387
rect 532 -390 538 -387
rect 544 -390 550 -387
rect 556 -390 562 -387
rect 568 -390 574 -387
rect 580 -390 586 -387
rect 592 -390 598 -387
rect 604 -390 610 -387
rect 616 -390 622 -387
rect 628 -390 634 -387
rect 640 -390 646 -387
rect 652 -390 658 -387
rect 664 -390 670 -387
rect 676 -390 682 -387
rect 688 -390 694 -387
rect 700 -390 706 -387
rect 712 -390 718 -387
rect 724 -390 730 -387
rect 736 -390 742 -387
rect 748 -390 754 -387
rect 760 -390 766 -387
rect 772 -390 778 -387
rect -606 -394 778 -390
<< polycontact >>
rect 16 130 20 134
rect 185 124 189 128
rect -15 114 -11 118
rect 26 1 30 5
rect 58 -1 62 3
rect 110 -1 114 3
rect 141 -1 145 3
rect 153 -9 157 -5
rect -593 -144 -589 -140
rect -581 -144 -577 -140
rect -569 -144 -565 -140
rect -557 -144 -553 -140
rect -545 -144 -541 -140
rect -533 -144 -529 -140
rect -521 -144 -517 -140
rect -509 -144 -505 -140
rect -497 -144 -493 -140
rect -485 -144 -481 -140
rect -473 -144 -469 -140
rect -461 -144 -457 -140
rect -449 -144 -445 -140
rect -437 -144 -433 -140
rect -425 -144 -421 -140
rect -413 -144 -409 -140
rect -401 -144 -397 -140
rect -389 -144 -385 -140
rect -377 -144 -373 -140
rect -365 -144 -361 -140
rect -353 -144 -349 -140
rect -341 -144 -337 -140
rect -329 -144 -325 -140
rect -317 -144 -313 -140
rect -305 -144 -301 -140
rect -293 -144 -289 -140
rect -281 -144 -277 -140
rect -269 -144 -265 -140
rect -257 -144 -253 -140
rect -245 -144 -241 -140
rect -233 -144 -229 -140
rect -221 -144 -217 -140
rect -209 -144 -205 -140
rect -197 -144 -193 -140
rect -185 -144 -181 -140
rect -173 -144 -169 -140
rect -161 -144 -157 -140
rect -149 -144 -145 -140
rect -137 -144 -133 -140
rect -125 -144 -121 -140
rect -113 -144 -109 -140
rect -101 -144 -97 -140
rect -89 -144 -85 -140
rect -77 -144 -73 -140
rect -65 -144 -61 -140
rect -53 -144 -49 -140
rect -41 -144 -37 -140
rect -29 -144 -25 -140
<< metal1 >>
rect -599 114 -19 117
rect -599 111 -595 114
rect -575 111 -571 114
rect -551 111 -547 114
rect -527 111 -523 114
rect -503 111 -499 114
rect -479 111 -475 114
rect -455 111 -451 114
rect -431 111 -427 114
rect -407 111 -403 114
rect -383 111 -379 114
rect -359 111 -355 114
rect -335 111 -331 114
rect -311 111 -307 114
rect -287 111 -283 114
rect -263 111 -259 114
rect -239 111 -235 114
rect -215 111 -211 114
rect -191 111 -187 114
rect -167 111 -163 114
rect -143 111 -139 114
rect -119 111 -115 114
rect -95 111 -91 114
rect -71 111 -67 114
rect -47 111 -43 114
rect -23 111 -19 114
rect -626 -132 -622 -130
rect 16 110 20 130
rect 46 122 50 126
rect 169 117 771 121
rect 191 114 195 117
rect 215 114 219 117
rect 239 114 243 117
rect 263 114 267 117
rect 287 114 291 117
rect 311 114 315 117
rect 335 114 339 117
rect 359 114 363 117
rect 383 114 387 117
rect 407 114 411 117
rect 431 114 435 117
rect 455 114 459 117
rect 479 114 483 117
rect 503 114 507 117
rect 527 114 531 117
rect 551 114 555 117
rect 575 114 579 117
rect 599 114 603 117
rect 623 114 627 117
rect 647 114 651 117
rect 671 114 675 117
rect 695 114 699 117
rect 719 114 723 117
rect 743 114 747 117
rect 767 114 771 117
rect 26 -1 30 1
rect 11 -5 30 -1
rect 58 -5 62 -1
rect 107 -5 114 -1
rect 141 -5 145 -1
rect 11 -10 15 -5
rect 103 -10 107 -5
rect 141 -9 153 -5
rect 165 -7 169 6
rect 46 -123 50 -119
rect -611 -132 -607 -129
rect -587 -132 -583 -129
rect -563 -132 -559 -129
rect -539 -132 -535 -129
rect -515 -132 -511 -129
rect -491 -132 -487 -129
rect -467 -132 -463 -129
rect -443 -132 -439 -129
rect -419 -132 -415 -129
rect -395 -132 -391 -129
rect -371 -132 -367 -129
rect -347 -132 -343 -129
rect -323 -132 -319 -129
rect -299 -132 -295 -129
rect -275 -132 -271 -129
rect -251 -132 -247 -129
rect -227 -132 -223 -129
rect -203 -132 -199 -129
rect -179 -132 -175 -129
rect -155 -132 -151 -129
rect -131 -132 -127 -129
rect -107 -132 -103 -129
rect -83 -132 -79 -129
rect -59 -132 -55 -129
rect -35 -132 -31 -129
rect -11 -132 -7 -129
rect -626 -136 -7 -132
rect 179 -129 183 -126
rect 203 -129 207 -126
rect 227 -129 231 -126
rect 251 -129 255 -126
rect 275 -129 279 -126
rect 299 -129 303 -126
rect 323 -129 327 -126
rect 347 -129 351 -126
rect 371 -129 375 -126
rect 395 -129 399 -126
rect 419 -129 423 -126
rect 443 -129 447 -126
rect 467 -129 471 -126
rect 491 -129 495 -126
rect 515 -129 519 -126
rect 539 -129 543 -126
rect 563 -129 567 -126
rect 587 -129 591 -126
rect 611 -129 615 -126
rect 635 -129 639 -126
rect 659 -129 663 -126
rect 683 -129 687 -126
rect 707 -129 711 -126
rect 731 -129 735 -126
rect 755 -129 759 -126
rect 779 -129 783 -126
rect 793 -129 797 -124
rect 179 -133 797 -129
rect 184 -136 778 -133
rect -599 -139 -19 -136
rect -620 -140 -19 -139
rect -620 -143 -593 -140
rect -599 -144 -593 -143
rect -589 -144 -581 -140
rect -577 -144 -569 -140
rect -565 -144 -557 -140
rect -553 -144 -545 -140
rect -541 -144 -533 -140
rect -529 -144 -521 -140
rect -517 -144 -509 -140
rect -505 -144 -497 -140
rect -493 -144 -485 -140
rect -481 -144 -473 -140
rect -469 -144 -461 -140
rect -457 -144 -449 -140
rect -445 -144 -437 -140
rect -433 -144 -425 -140
rect -421 -144 -413 -140
rect -409 -144 -401 -140
rect -397 -144 -389 -140
rect -385 -144 -377 -140
rect -373 -144 -365 -140
rect -361 -144 -353 -140
rect -349 -144 -341 -140
rect -337 -144 -329 -140
rect -325 -144 -317 -140
rect -313 -144 -305 -140
rect -301 -144 -293 -140
rect -289 -144 -281 -140
rect -277 -144 -269 -140
rect -265 -144 -257 -140
rect -253 -144 -245 -140
rect -241 -144 -233 -140
rect -229 -144 -221 -140
rect -217 -144 -209 -140
rect -205 -144 -197 -140
rect -193 -144 -185 -140
rect -181 -144 -173 -140
rect -169 -144 -161 -140
rect -157 -144 -149 -140
rect -145 -144 -137 -140
rect -133 -144 -125 -140
rect -121 -144 -113 -140
rect -109 -144 -101 -140
rect -97 -144 -89 -140
rect -85 -144 -77 -140
rect -73 -144 -65 -140
rect -61 -144 -53 -140
rect -49 -144 -41 -140
rect -37 -144 -29 -140
rect -25 -144 -19 -140
rect -599 -147 -595 -144
rect -575 -147 -571 -144
rect -551 -147 -547 -144
rect -527 -147 -523 -144
rect -503 -147 -499 -144
rect -479 -147 -475 -144
rect -455 -147 -451 -144
rect -431 -147 -427 -144
rect -407 -147 -403 -144
rect -383 -147 -379 -144
rect -359 -147 -355 -144
rect -335 -147 -331 -144
rect -311 -147 -307 -144
rect -287 -147 -283 -144
rect -263 -147 -259 -144
rect -239 -147 -235 -144
rect -215 -147 -211 -144
rect -191 -147 -187 -144
rect -167 -147 -163 -144
rect -143 -147 -139 -144
rect -119 -147 -115 -144
rect -95 -147 -91 -144
rect -71 -147 -67 -144
rect -47 -147 -43 -144
rect -23 -147 -19 -144
rect 191 -144 778 -136
rect 191 -147 195 -144
rect 215 -147 219 -144
rect 239 -147 243 -144
rect 263 -147 267 -144
rect 287 -147 291 -144
rect 311 -147 315 -144
rect 335 -147 339 -144
rect 359 -147 363 -144
rect 383 -147 387 -144
rect 407 -147 411 -144
rect 431 -147 435 -144
rect 455 -147 459 -144
rect 479 -147 483 -144
rect 503 -147 507 -144
rect 527 -147 531 -144
rect 551 -147 555 -144
rect 575 -147 579 -144
rect 599 -147 603 -144
rect 623 -147 627 -144
rect 647 -147 651 -144
rect 671 -147 675 -144
rect 695 -147 699 -144
rect 719 -147 723 -144
rect 743 -147 747 -144
rect 767 -147 771 -144
rect -611 -390 -607 -387
rect -587 -390 -583 -387
rect -563 -390 -559 -387
rect -539 -390 -535 -387
rect -515 -390 -511 -387
rect -491 -390 -487 -387
rect -467 -390 -463 -387
rect -443 -390 -439 -387
rect -419 -390 -415 -387
rect -395 -390 -391 -387
rect -371 -390 -367 -387
rect -347 -390 -343 -387
rect -323 -390 -319 -387
rect -299 -390 -295 -387
rect -275 -390 -271 -387
rect -251 -390 -247 -387
rect -227 -390 -223 -387
rect -203 -390 -199 -387
rect -179 -390 -175 -387
rect -155 -390 -151 -387
rect -131 -390 -127 -387
rect -107 -390 -103 -387
rect -83 -390 -79 -387
rect -59 -390 -55 -387
rect -35 -390 -31 -387
rect -11 -390 -7 -387
rect 5 -268 9 -264
rect 5 -390 9 -383
rect -611 -394 9 -390
rect 165 -269 169 -265
rect 165 -390 169 -383
rect 179 -390 183 -387
rect 203 -390 207 -387
rect 227 -390 231 -387
rect 251 -390 255 -387
rect 275 -390 279 -387
rect 299 -390 303 -387
rect 323 -390 327 -387
rect 347 -390 351 -387
rect 371 -390 375 -387
rect 395 -390 399 -387
rect 419 -390 423 -387
rect 443 -390 447 -387
rect 467 -390 471 -387
rect 491 -390 495 -387
rect 515 -390 519 -387
rect 539 -390 543 -387
rect 563 -390 567 -387
rect 587 -390 591 -387
rect 611 -390 615 -387
rect 635 -390 639 -387
rect 659 -390 663 -387
rect 683 -390 687 -387
rect 707 -390 711 -387
rect 731 -390 735 -387
rect 755 -390 759 -387
rect 779 -390 783 -387
rect 165 -394 783 -390
<< m2contact >>
rect 131 251 135 255
rect -11 114 -7 118
rect -19 -22 -15 -18
rect 185 128 189 132
rect 122 122 126 126
rect 15 106 19 110
rect 37 6 41 10
rect 103 -5 107 -1
rect 1 -22 5 -18
rect 122 -153 126 -149
<< metal2 >>
rect 131 132 135 251
rect 131 128 185 132
rect -7 114 41 118
rect 15 -1 19 106
rect 37 10 41 114
rect 15 -5 103 -1
rect -15 -22 1 -18
rect 122 -149 126 122
use amp  amp_0
timestamp 1418875346
transform 1 0 95 0 1 135
box -95 -135 77 126
use bias  bias_0
timestamp 1418768461
transform 1 0 -11 0 1 -106
box 13 -282 183 102
<< labels >>
rlabel metal1 -611 -394 -607 -390 1 Gnd
rlabel space 76 13 80 17 1 V-p
rlabel space 33 6 37 10 1 V-fb
rlabel space 135 6 139 10 1 V-fb
rlabel space 92 13 96 17 1 V-n
rlabel space 76 244 80 248 1 V+p
rlabel space 92 244 96 248 1 V+n
rlabel space 33 251 37 255 1 V+fb
rlabel space 135 251 139 255 1 V+fb
rlabel metal1 -599 -142 -595 -138 1 Vout_not
<< end >>
