magic
tech scmos
timestamp 1418882595
<< nwell >>
rect 1556 1421 1560 1425
<< polysilicon >>
rect 1556 1421 1560 1424
<< polycontact >>
rect 1556 1424 1560 1428
<< m2contact >>
rect 738 1471 742 1475
rect 1552 1424 1556 1428
<< metal2 >>
rect 1544 4511 1558 4527
rect 641 4443 656 4448
rect 653 4433 656 4443
rect 1071 4443 1085 4511
rect 4389 4448 4403 4492
rect 1071 4439 1072 4443
rect 1080 4439 1085 4443
rect 4365 4434 4403 4448
rect 641 4336 656 4433
rect 641 4313 662 4336
rect 642 1455 662 4313
rect 4365 1530 4370 4434
rect 4365 1522 4370 1523
rect 4391 4403 4470 4404
rect 4391 4389 4509 4403
rect 4391 4388 4470 4389
rect 4391 1515 4398 4388
rect 4401 3914 4499 3930
rect 4391 1510 4392 1515
rect 4397 1510 4398 1515
rect 4391 1509 4398 1510
rect 4402 1506 4407 3914
rect 4402 1500 4407 1501
rect 4411 3440 4491 3456
rect 4411 1497 4416 3440
rect 4420 2966 4500 2982
rect 4411 1492 4412 1497
rect 4411 1491 4416 1492
rect 4420 1487 4425 2966
rect 4424 1482 4425 1487
rect 4420 1481 4425 1482
rect 738 1475 742 1476
rect 642 1451 1550 1455
rect 645 1449 722 1451
rect 1446 1434 1453 1439
rect 1446 1432 1449 1434
rect 1450 1410 1454 1417
rect 1476 1415 1479 1420
rect 4398 732 4399 739
rect 2965 723 2978 724
rect 2965 717 2967 723
rect 2965 638 2978 717
rect 4392 710 4399 732
rect 3441 709 3454 710
rect 3441 702 3443 709
rect 3453 702 3454 709
rect 2964 517 2980 638
rect 3441 633 3454 702
rect 3918 641 3928 688
rect 4392 649 4399 701
rect 2965 506 2980 517
rect 2964 485 2980 506
rect 3439 480 3455 633
rect 3914 488 3930 641
rect 4388 496 4404 649
<< m3contact >>
rect 641 4433 653 4443
rect 1072 4434 1080 4443
rect 4364 1523 4370 1530
rect 4392 1510 4397 1515
rect 4402 1501 4407 1506
rect 4412 1492 4417 1497
rect 4419 1482 4424 1487
rect 738 1476 743 1481
rect 1470 1440 1475 1445
rect 1449 1429 1454 1434
rect 1460 1423 1465 1429
rect 1479 1415 1484 1420
rect 1396 1372 1401 1377
rect 1396 1348 1401 1353
rect 1396 1324 1401 1329
rect 1396 1300 1401 1305
rect 4391 732 4398 739
rect 2967 717 2978 723
rect 3443 702 3453 709
rect 3916 688 3928 694
<< metal3 >>
rect 638 4443 1087 4447
rect 638 4433 641 4443
rect 653 4434 1072 4443
rect 1080 4434 1087 4443
rect 653 4433 1087 4434
rect 638 4432 1087 4433
rect 1069 4431 1087 4432
rect 4363 1530 4371 1531
rect 4363 1529 4364 1530
rect 738 1523 4364 1529
rect 4370 1523 4371 1530
rect 739 1482 744 1523
rect 4363 1522 4371 1523
rect 4391 1515 4398 1516
rect 737 1481 744 1482
rect 737 1476 738 1481
rect 743 1476 744 1481
rect 737 1475 744 1476
rect 1397 1510 4392 1515
rect 4397 1510 4398 1515
rect 1397 1509 4398 1510
rect 1397 1378 1402 1509
rect 4401 1506 4408 1507
rect 1395 1377 1402 1378
rect 1395 1372 1396 1377
rect 1401 1372 1402 1377
rect 1395 1371 1402 1372
rect 1405 1501 4402 1506
rect 4407 1501 4408 1506
rect 1405 1500 4408 1501
rect 1395 1353 1402 1354
rect 1395 1348 1396 1353
rect 1401 1352 1402 1353
rect 1405 1352 1410 1500
rect 4411 1497 4418 1498
rect 1401 1348 1410 1352
rect 1395 1347 1410 1348
rect 1413 1492 4412 1497
rect 4417 1492 4418 1497
rect 1413 1491 4418 1492
rect 1395 1329 1402 1330
rect 1395 1324 1396 1329
rect 1401 1328 1402 1329
rect 1413 1328 1418 1491
rect 1401 1324 1418 1328
rect 1395 1323 1418 1324
rect 1421 1487 4425 1488
rect 1421 1482 4419 1487
rect 4424 1482 4425 1487
rect 1395 1305 1402 1306
rect 1395 1300 1396 1305
rect 1401 1304 1402 1305
rect 1421 1304 1426 1482
rect 4418 1481 4425 1482
rect 1469 1445 1476 1446
rect 1469 1440 1470 1445
rect 1475 1440 1476 1445
rect 1469 1439 1476 1440
rect 1448 1434 1455 1435
rect 1448 1429 1449 1434
rect 1454 1429 1455 1434
rect 1448 1413 1455 1429
rect 1459 1429 1466 1430
rect 1459 1423 1460 1429
rect 1465 1423 1466 1429
rect 1459 1422 1466 1423
rect 1401 1300 1434 1304
rect 1395 1299 1434 1300
rect 1450 711 1455 1413
rect 1449 696 1455 711
rect 1461 710 1466 1422
rect 1469 724 1474 1439
rect 1478 1420 1485 1421
rect 1477 1415 1479 1420
rect 1484 1415 1485 1420
rect 1477 1414 1485 1415
rect 1477 1413 1484 1414
rect 1477 740 1482 1413
rect 1477 739 4447 740
rect 1477 732 4391 739
rect 4398 732 4447 739
rect 1477 731 4447 732
rect 1469 723 4445 724
rect 1469 717 2967 723
rect 2978 717 4445 723
rect 1469 715 4445 717
rect 1461 709 4437 710
rect 1461 702 3443 709
rect 3453 702 4437 709
rect 1461 701 4437 702
rect 1449 694 4427 696
rect 1449 688 3916 694
rect 3928 688 4427 694
rect 1449 687 4427 688
use barepad  barepad_1
timestamp 1259953556
transform -1 0 841 0 -1 5000
box -2 0 476 513
use inpad  inpad_1
timestamp 1259953556
transform -1 0 1315 0 -1 5000
box -2 0 476 513
use inpad  inpad_0
timestamp 1259953556
transform -1 0 1789 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_3
timestamp 1259953556
transform -1 0 2263 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_6
timestamp 1259953556
transform -1 0 2737 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_5
timestamp 1259953556
transform -1 0 3211 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_4
timestamp 1259953556
transform -1 0 3685 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_3
timestamp 1259953556
transform -1 0 4159 0 -1 5000
box -2 0 476 513
use barepad  barepad_0
timestamp 1259953556
transform -1 0 4633 0 -1 5000
box -2 0 476 513
use padframe_top  padframe_top_0
timestamp 1259953556
transform 1 0 0 0 1 4487
box 0 0 5000 513
use barepad  barepad_2
timestamp 1259953556
transform 0 1 0 -1 0 4633
box -2 0 476 513
use inorpad  inorpad_7
timestamp 1259953556
transform 0 1 0 -1 0 4159
box -2 0 476 513
use inorpad  inorpad_8
timestamp 1259953556
transform 0 1 0 -1 0 3685
box -2 0 476 513
use inorpad  inorpad_9
timestamp 1259953556
transform 0 1 0 -1 0 3211
box -2 0 476 513
use inorpad  inorpad_10
timestamp 1259953556
transform 0 1 0 -1 0 2737
box -2 0 476 513
use inpad  inpad_2
timestamp 1259953556
transform 0 1 0 -1 0 2263
box -2 0 476 513
use inorpad  inorpad_17
timestamp 1259953556
transform 0 -1 5000 1 0 4159
box -2 0 476 513
use inorpad  inorpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 3685
box -2 0 476 513
use inorpad  inorpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 3211
box -2 0 476 513
use inorpad  inorpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 2737
box -2 0 476 513
use blankpad  blankpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 2263
box -2 0 476 513
use blankpad  blankpad_7
timestamp 1259953556
transform 0 -1 5000 1 0 1789
box -2 0 476 513
use inpad  inpad_3
timestamp 1259953556
transform 0 1 0 -1 0 1789
box -2 0 476 513
use inpad  inpad_4
timestamp 1259953556
transform 0 1 0 -1 0 1315
box -2 0 476 513
use top-level  top-level_0
timestamp 1418882011
transform 1 0 705 0 1 772
box 0 0 1733 711
use top-level  top-level_1
timestamp 1418882011
transform 1 0 2594 0 1 771
box 0 0 1733 711
use blankpad  blankpad_8
timestamp 1259953556
transform 0 -1 5000 1 0 1315
box -2 0 476 513
use blankpad  blankpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 841
box -2 0 476 513
use padframe_left  padframe_left_0
timestamp 1259953556
transform 1 0 0 0 1 367
box 2 2 513 4264
use iopad  iopad_0
timestamp 1259953556
transform 0 1 0 -1 0 841
box -2 0 476 513
use iopad  iopad_1
timestamp 1259953556
transform 1 0 367 0 1 0
box -2 0 476 513
use inorpad  inorpad_11
timestamp 1259953556
transform 1 0 841 0 1 0
box -2 0 476 513
use inorpad  inorpad_12
timestamp 1259953556
transform 1 0 1315 0 1 0
box -2 0 476 513
use iopad  iopad_2
timestamp 1259953556
transform 1 0 1789 0 1 0
box -2 0 476 513
use iopad  iopad_3
timestamp 1259953556
transform 1 0 2263 0 1 0
box -2 0 476 513
use inorpad  inorpad_13
timestamp 1259953556
transform 1 0 2737 0 1 0
box -2 0 476 513
use inorpad  inorpad_14
timestamp 1259953556
transform 1 0 3211 0 1 0
box -2 0 476 513
use inorpad  inorpad_15
timestamp 1259953556
transform 1 0 3685 0 1 0
box -2 0 476 513
use padframe_right  padframe_right_0
timestamp 1259953556
transform 1 0 4487 0 1 367
box 0 2 511 4264
use blankpad  blankpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 367
box -2 0 476 513
use inorpad  inorpad_16
timestamp 1259953556
transform 1 0 4159 0 1 0
box -2 0 476 513
use padframe_bottom  padframe_bottom_0
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 5000 513
<< labels >>
rlabel space 1396 1415 1402 1418 1 x1
rlabel space 1404 1415 1410 1418 1 x2
rlabel space 1412 1415 1418 1418 1 x3
rlabel space 1420 1415 1426 1418 1 x4
<< end >>
