magic
tech scmos
timestamp 1418869571
<< nwell >>
rect 2429 632 2453 648
rect 2485 632 2509 648
rect 2429 627 2462 632
rect 766 603 770 607
rect 766 599 769 600
rect 766 579 770 583
rect 518 511 562 514
rect 636 511 670 514
rect 2418 511 2462 627
rect 2536 622 2570 627
rect 2536 523 2612 622
rect 2664 523 2681 622
rect 2536 511 2570 523
rect 2063 390 2681 511
rect 2724 390 2767 655
rect 2810 514 2853 655
rect 2810 390 3471 514
rect 2063 258 3471 390
<< pwell >>
rect 2453 632 2485 648
rect 753 618 756 619
rect 761 613 762 614
rect 759 612 762 613
rect 759 611 761 612
rect 760 608 761 611
rect 752 604 753 607
rect 760 597 763 608
rect 2381 514 2412 627
rect 2472 627 2491 632
rect 2472 514 2536 627
rect 2612 523 2664 622
rect 2681 390 2724 655
rect 2767 390 2810 655
rect 2063 6 3471 258
rect 2063 1 2683 6
rect 2846 5 3471 6
rect 2846 4 2860 5
<< electrode >>
rect 1932 695 1940 700
rect 2340 695 2350 700
rect 2550 695 2560 700
rect 2610 695 2620 700
rect 2720 695 2730 700
rect 2780 695 2791 700
rect 3583 695 3591 700
rect 1932 694 1938 695
rect 2342 694 2348 695
rect 2552 694 2558 695
rect 2612 694 2618 695
rect 2722 694 2728 695
rect 2782 694 2788 695
rect 3585 694 3591 695
rect 2772 118 2778 125
rect 2772 87 2778 94
<< electrodecontact >>
rect 1933 695 1937 699
rect 2343 695 2347 699
rect 2553 695 2557 699
rect 2613 695 2617 699
rect 2723 695 2727 699
rect 2783 695 2787 699
rect 3586 695 3590 699
rect 1686 268 1690 420
rect 2055 264 2059 416
rect 3474 270 3478 420
rect 3586 268 3590 420
rect 2773 120 2777 124
rect 2773 88 2777 92
<< electrodecap >>
rect 1905 262 2061 418
rect 3472 266 3628 422
<< ntransistor >>
rect 2173 684 2338 686
rect 2383 684 2548 686
rect 2796 684 2961 686
rect 2971 684 3136 686
rect 2464 638 2466 642
rect 2472 638 2474 642
rect 2399 612 2401 616
rect 2392 607 2394 611
rect 2483 615 2491 619
rect 2494 615 2502 619
rect 2520 612 2522 616
rect 2399 601 2401 605
rect 2483 607 2491 611
rect 2494 607 2502 611
rect 2520 601 2522 605
rect 2399 585 2401 589
rect 2392 580 2394 584
rect 2483 588 2491 592
rect 2494 588 2502 592
rect 2520 585 2522 589
rect 2399 574 2401 578
rect 2483 580 2491 584
rect 2494 580 2502 584
rect 2626 612 2628 616
rect 2633 606 2635 610
rect 2654 608 2658 610
rect 2626 601 2628 605
rect 2520 574 2522 578
rect 2626 588 2628 592
rect 2399 558 2401 562
rect 2392 553 2394 557
rect 2483 561 2491 565
rect 2494 561 2502 565
rect 2520 558 2522 562
rect 2399 547 2401 551
rect 2483 553 2491 557
rect 2494 553 2502 557
rect 2633 582 2635 586
rect 2654 584 2658 586
rect 2626 577 2628 581
rect 2626 564 2628 568
rect 2520 547 2522 551
rect 2399 531 2401 535
rect 2392 526 2394 530
rect 2483 534 2491 538
rect 2494 534 2502 538
rect 2520 531 2522 535
rect 2399 520 2401 524
rect 2483 526 2491 530
rect 2494 526 2502 530
rect 2633 558 2635 562
rect 2654 560 2658 562
rect 2626 553 2628 557
rect 2626 540 2628 544
rect 2520 520 2522 524
rect 2633 534 2635 538
rect 2654 536 2658 538
rect 2626 529 2628 533
rect 2695 529 2701 649
rect 2707 529 2713 649
rect 2778 529 2784 649
rect 2695 400 2701 520
rect 2707 400 2713 520
rect 2778 400 2784 520
rect 2790 400 2796 520
rect 2075 7 2081 247
rect 2087 7 2093 247
rect 2099 7 2105 247
rect 2111 7 2117 247
rect 2123 7 2129 247
rect 2135 7 2141 247
rect 2147 7 2153 247
rect 2159 7 2165 247
rect 2171 7 2177 247
rect 2183 7 2189 247
rect 2195 7 2201 247
rect 2207 7 2213 247
rect 2219 7 2225 247
rect 2231 7 2237 247
rect 2243 7 2249 247
rect 2255 7 2261 247
rect 2267 7 2273 247
rect 2279 7 2285 247
rect 2291 7 2297 247
rect 2303 7 2309 247
rect 2315 7 2321 247
rect 2327 7 2333 247
rect 2339 7 2345 247
rect 2351 7 2357 247
rect 2363 7 2369 247
rect 2375 7 2381 247
rect 2387 7 2393 247
rect 2399 7 2405 247
rect 2411 7 2417 247
rect 2423 7 2429 247
rect 2435 7 2441 247
rect 2447 7 2453 247
rect 2459 7 2465 247
rect 2471 7 2477 247
rect 2483 7 2489 247
rect 2495 7 2501 247
rect 2507 7 2513 247
rect 2519 7 2525 247
rect 2531 7 2537 247
rect 2543 7 2549 247
rect 2555 7 2561 247
rect 2567 7 2573 247
rect 2579 7 2585 247
rect 2591 7 2597 247
rect 2603 7 2609 247
rect 2615 7 2621 247
rect 2627 7 2633 247
rect 2639 7 2645 247
rect 2651 7 2657 247
rect 2663 7 2669 247
rect 2697 132 2703 252
rect 2709 132 2715 252
rect 2721 132 2727 252
rect 2733 132 2739 252
rect 2753 12 2759 252
rect 2777 132 2783 252
rect 2797 132 2803 252
rect 2809 132 2815 252
rect 2821 132 2827 252
rect 2833 132 2839 252
rect 2865 11 2871 251
rect 2877 11 2883 251
rect 2889 11 2895 251
rect 2901 11 2907 251
rect 2913 11 2919 251
rect 2925 11 2931 251
rect 2937 11 2943 251
rect 2949 11 2955 251
rect 2961 11 2967 251
rect 2973 11 2979 251
rect 2985 11 2991 251
rect 2997 11 3003 251
rect 3009 11 3015 251
rect 3021 11 3027 251
rect 3033 11 3039 251
rect 3045 11 3051 251
rect 3057 11 3063 251
rect 3069 11 3075 251
rect 3081 11 3087 251
rect 3093 11 3099 251
rect 3105 11 3111 251
rect 3117 11 3123 251
rect 3129 11 3135 251
rect 3141 11 3147 251
rect 3153 11 3159 251
rect 3165 11 3171 251
rect 3177 11 3183 251
rect 3189 11 3195 251
rect 3201 11 3207 251
rect 3213 11 3219 251
rect 3225 11 3231 251
rect 3237 11 3243 251
rect 3249 11 3255 251
rect 3261 11 3267 251
rect 3273 11 3279 251
rect 3285 11 3291 251
rect 3297 11 3303 251
rect 3309 11 3315 251
rect 3321 11 3327 251
rect 3333 11 3339 251
rect 3345 11 3351 251
rect 3357 11 3363 251
rect 3369 11 3375 251
rect 3381 11 3387 251
rect 3393 11 3399 251
rect 3405 11 3411 251
rect 3417 11 3423 251
rect 3429 11 3435 251
rect 3441 11 3447 251
rect 3453 11 3459 251
<< ptransistor >>
rect 2440 638 2442 642
rect 2496 638 2498 642
rect 2429 612 2431 616
rect 2449 615 2451 619
rect 2449 607 2451 611
rect 2550 612 2552 616
rect 2429 601 2431 605
rect 2576 612 2578 616
rect 2596 612 2598 616
rect 2557 606 2559 610
rect 2550 601 2552 605
rect 2429 585 2431 589
rect 2449 588 2451 592
rect 2449 580 2451 584
rect 2550 585 2552 589
rect 2429 574 2431 578
rect 2576 601 2578 605
rect 2596 601 2598 605
rect 2670 608 2674 610
rect 2576 588 2578 592
rect 2596 588 2598 592
rect 2557 579 2559 583
rect 2550 574 2552 578
rect 2429 558 2431 562
rect 2449 561 2451 565
rect 2449 553 2451 557
rect 2550 558 2552 562
rect 2429 547 2431 551
rect 2576 577 2578 581
rect 2596 577 2598 581
rect 2670 584 2674 586
rect 2576 564 2578 568
rect 2596 564 2598 568
rect 2557 552 2559 556
rect 2576 553 2578 557
rect 2596 553 2598 557
rect 2550 547 2552 551
rect 2429 531 2431 535
rect 2449 534 2451 538
rect 2449 526 2451 530
rect 2550 531 2552 535
rect 2429 520 2431 524
rect 2670 560 2674 562
rect 2576 540 2578 544
rect 2596 540 2598 544
rect 2576 529 2578 533
rect 2596 529 2598 533
rect 2557 525 2559 529
rect 2550 520 2552 524
rect 2670 536 2674 538
rect 2750 529 2756 649
rect 2821 529 2827 649
rect 2833 529 2839 649
rect 2075 265 2081 505
rect 2087 265 2093 505
rect 2099 265 2105 505
rect 2111 265 2117 505
rect 2123 265 2129 505
rect 2135 265 2141 505
rect 2147 265 2153 505
rect 2159 265 2165 505
rect 2171 265 2177 505
rect 2183 265 2189 505
rect 2195 265 2201 505
rect 2207 265 2213 505
rect 2219 265 2225 505
rect 2231 265 2237 505
rect 2243 265 2249 505
rect 2255 265 2261 505
rect 2267 265 2273 505
rect 2279 265 2285 505
rect 2291 265 2297 505
rect 2303 265 2309 505
rect 2315 265 2321 505
rect 2327 265 2333 505
rect 2339 265 2345 505
rect 2351 265 2357 505
rect 2363 265 2369 505
rect 2375 265 2381 505
rect 2387 265 2393 505
rect 2399 265 2405 505
rect 2411 265 2417 505
rect 2423 265 2429 505
rect 2435 265 2441 505
rect 2447 265 2453 505
rect 2459 265 2465 505
rect 2471 265 2477 505
rect 2483 265 2489 505
rect 2495 265 2501 505
rect 2507 265 2513 505
rect 2519 265 2525 505
rect 2531 265 2537 505
rect 2543 265 2549 505
rect 2555 265 2561 505
rect 2567 265 2573 505
rect 2579 265 2585 505
rect 2591 265 2597 505
rect 2603 265 2609 505
rect 2615 265 2621 505
rect 2627 265 2633 505
rect 2639 265 2645 505
rect 2651 265 2657 505
rect 2663 265 2669 505
rect 2738 400 2744 520
rect 2750 400 2756 520
rect 2821 400 2827 520
rect 2833 400 2839 520
rect 2697 264 2703 384
rect 2709 264 2715 384
rect 2721 264 2727 384
rect 2733 264 2739 384
rect 2753 264 2759 384
rect 2777 264 2783 384
rect 2797 264 2803 384
rect 2809 264 2815 384
rect 2821 264 2827 384
rect 2833 264 2839 384
rect 2865 268 2871 508
rect 2877 268 2883 508
rect 2889 268 2895 508
rect 2901 268 2907 508
rect 2913 268 2919 508
rect 2925 268 2931 508
rect 2937 268 2943 508
rect 2949 268 2955 508
rect 2961 268 2967 508
rect 2973 268 2979 508
rect 2985 268 2991 508
rect 2997 268 3003 508
rect 3009 268 3015 508
rect 3021 268 3027 508
rect 3033 268 3039 508
rect 3045 268 3051 508
rect 3057 268 3063 508
rect 3069 268 3075 508
rect 3081 268 3087 508
rect 3093 268 3099 508
rect 3105 268 3111 508
rect 3117 268 3123 508
rect 3129 268 3135 508
rect 3141 268 3147 508
rect 3153 268 3159 508
rect 3165 268 3171 508
rect 3177 268 3183 508
rect 3189 268 3195 508
rect 3201 268 3207 508
rect 3213 268 3219 508
rect 3225 268 3231 508
rect 3237 268 3243 508
rect 3249 268 3255 508
rect 3261 268 3267 508
rect 3273 268 3279 508
rect 3285 268 3291 508
rect 3297 268 3303 508
rect 3309 268 3315 508
rect 3321 268 3327 508
rect 3333 268 3339 508
rect 3345 268 3351 508
rect 3357 268 3363 508
rect 3369 268 3375 508
rect 3381 268 3387 508
rect 3393 268 3399 508
rect 3405 268 3411 508
rect 3417 268 3423 508
rect 3429 268 3435 508
rect 3441 268 3447 508
rect 3453 268 3459 508
<< ndiffusion >>
rect 2177 687 2338 689
rect 2173 686 2338 687
rect 2387 687 2548 689
rect 2383 686 2548 687
rect 2800 687 2961 689
rect 2796 686 2961 687
rect 2975 687 3136 689
rect 2971 686 3136 687
rect 2173 683 2338 684
rect 2173 681 2334 683
rect 2383 683 2548 684
rect 2383 681 2544 683
rect 2796 683 2961 684
rect 2971 683 3136 684
rect 2796 681 2802 683
rect 2806 681 3136 683
rect 2958 680 2974 681
rect 2463 638 2464 642
rect 2466 638 2467 642
rect 2471 638 2472 642
rect 2474 638 2475 642
rect 2388 611 2391 612
rect 2395 612 2399 616
rect 2401 612 2402 616
rect 2395 611 2398 612
rect 2388 607 2392 611
rect 2394 607 2398 611
rect 2482 615 2483 619
rect 2491 615 2494 619
rect 2502 615 2503 619
rect 2388 605 2391 607
rect 2388 584 2391 585
rect 2395 605 2398 607
rect 2519 612 2520 616
rect 2522 612 2523 616
rect 2395 601 2399 605
rect 2401 601 2402 605
rect 2482 607 2483 611
rect 2491 607 2494 611
rect 2502 607 2503 611
rect 2519 601 2520 605
rect 2522 601 2523 605
rect 2395 585 2399 589
rect 2401 585 2402 589
rect 2395 584 2398 585
rect 2388 580 2392 584
rect 2394 580 2398 584
rect 2482 588 2483 592
rect 2491 588 2494 592
rect 2502 588 2503 592
rect 2388 578 2391 580
rect 2388 557 2391 558
rect 2395 578 2398 580
rect 2519 585 2520 589
rect 2522 585 2523 589
rect 2395 574 2399 578
rect 2401 574 2402 578
rect 2482 580 2483 584
rect 2491 580 2494 584
rect 2502 580 2503 584
rect 2625 612 2626 616
rect 2628 612 2632 616
rect 2629 610 2632 612
rect 2636 610 2639 612
rect 2629 606 2633 610
rect 2635 606 2639 610
rect 2654 610 2658 611
rect 2629 605 2632 606
rect 2625 601 2626 605
rect 2628 601 2632 605
rect 2519 574 2520 578
rect 2522 574 2523 578
rect 2625 588 2626 592
rect 2628 588 2632 592
rect 2629 586 2632 588
rect 2636 605 2639 606
rect 2654 607 2658 608
rect 2636 586 2639 588
rect 2395 558 2399 562
rect 2401 558 2402 562
rect 2395 557 2398 558
rect 2388 553 2392 557
rect 2394 553 2398 557
rect 2482 561 2483 565
rect 2491 561 2494 565
rect 2502 561 2503 565
rect 2388 551 2391 553
rect 2388 530 2391 531
rect 2395 551 2398 553
rect 2519 558 2520 562
rect 2522 558 2523 562
rect 2395 547 2399 551
rect 2401 547 2402 551
rect 2482 553 2483 557
rect 2491 553 2494 557
rect 2502 553 2503 557
rect 2629 582 2633 586
rect 2635 582 2639 586
rect 2654 586 2658 587
rect 2629 581 2632 582
rect 2625 577 2626 581
rect 2628 577 2632 581
rect 2625 564 2626 568
rect 2628 564 2632 568
rect 2629 562 2632 564
rect 2636 581 2639 582
rect 2654 583 2658 584
rect 2636 562 2639 564
rect 2519 547 2520 551
rect 2522 547 2523 551
rect 2395 531 2399 535
rect 2401 531 2402 535
rect 2395 530 2398 531
rect 2388 526 2392 530
rect 2394 526 2398 530
rect 2482 534 2483 538
rect 2491 534 2494 538
rect 2502 534 2503 538
rect 2388 524 2391 526
rect 2395 524 2398 526
rect 2519 531 2520 535
rect 2522 531 2523 535
rect 2395 520 2399 524
rect 2401 520 2402 524
rect 2482 526 2483 530
rect 2491 526 2494 530
rect 2502 526 2503 530
rect 2629 558 2633 562
rect 2635 558 2639 562
rect 2654 562 2658 563
rect 2629 557 2632 558
rect 2625 553 2626 557
rect 2628 553 2632 557
rect 2625 540 2626 544
rect 2628 540 2632 544
rect 2629 538 2632 540
rect 2636 557 2639 558
rect 2654 559 2658 560
rect 2636 538 2639 540
rect 2519 520 2520 524
rect 2522 520 2523 524
rect 2629 534 2633 538
rect 2635 534 2639 538
rect 2654 538 2658 539
rect 2629 533 2632 534
rect 2625 529 2626 533
rect 2628 529 2632 533
rect 2636 533 2639 534
rect 2654 535 2658 536
rect 2692 533 2695 649
rect 2694 529 2695 533
rect 2701 642 2707 649
rect 2701 638 2702 642
rect 2706 638 2707 642
rect 2701 529 2707 638
rect 2713 645 2714 649
rect 2713 529 2716 645
rect 2775 642 2778 649
rect 2777 638 2778 642
rect 2775 529 2778 638
rect 2784 533 2787 649
rect 2784 529 2785 533
rect 2694 516 2695 520
rect 2692 400 2695 516
rect 2701 411 2707 520
rect 2701 407 2702 411
rect 2706 407 2707 411
rect 2701 400 2707 407
rect 2713 404 2716 520
rect 2713 400 2714 404
rect 2775 411 2778 520
rect 2777 407 2778 411
rect 2775 400 2778 407
rect 2784 516 2785 520
rect 2789 516 2790 520
rect 2784 400 2790 516
rect 2796 516 2797 520
rect 2796 400 2799 516
rect 2694 250 2697 252
rect 2069 7 2070 247
rect 2074 7 2075 247
rect 2081 7 2082 247
rect 2086 7 2087 247
rect 2093 7 2094 247
rect 2098 7 2099 247
rect 2105 7 2106 247
rect 2110 7 2111 247
rect 2117 7 2118 247
rect 2122 7 2123 247
rect 2129 7 2130 247
rect 2134 7 2135 247
rect 2141 7 2142 247
rect 2146 7 2147 247
rect 2153 7 2154 247
rect 2158 7 2159 247
rect 2165 7 2166 247
rect 2170 7 2171 247
rect 2177 7 2178 247
rect 2182 7 2183 247
rect 2189 7 2190 247
rect 2194 7 2195 247
rect 2201 7 2202 247
rect 2206 7 2207 247
rect 2213 7 2214 247
rect 2218 7 2219 247
rect 2225 7 2226 247
rect 2230 7 2231 247
rect 2237 7 2238 247
rect 2242 7 2243 247
rect 2249 7 2250 247
rect 2254 7 2255 247
rect 2261 7 2262 247
rect 2266 7 2267 247
rect 2273 7 2274 247
rect 2278 7 2279 247
rect 2285 7 2286 247
rect 2290 7 2291 247
rect 2297 7 2298 247
rect 2302 7 2303 247
rect 2309 7 2310 247
rect 2314 7 2315 247
rect 2321 7 2322 247
rect 2326 7 2327 247
rect 2333 7 2334 247
rect 2338 7 2339 247
rect 2345 7 2346 247
rect 2350 7 2351 247
rect 2357 7 2358 247
rect 2362 7 2363 247
rect 2369 7 2370 247
rect 2374 7 2375 247
rect 2381 7 2382 247
rect 2386 7 2387 247
rect 2393 7 2394 247
rect 2398 7 2399 247
rect 2405 7 2406 247
rect 2410 7 2411 247
rect 2417 7 2418 247
rect 2422 7 2423 247
rect 2429 7 2430 247
rect 2434 7 2435 247
rect 2441 7 2442 247
rect 2446 7 2447 247
rect 2453 7 2454 247
rect 2458 7 2459 247
rect 2465 7 2466 247
rect 2470 7 2471 247
rect 2477 7 2478 247
rect 2482 7 2483 247
rect 2489 7 2490 247
rect 2494 7 2495 247
rect 2501 7 2502 247
rect 2506 7 2507 247
rect 2513 7 2514 247
rect 2518 7 2519 247
rect 2525 7 2526 247
rect 2530 7 2531 247
rect 2537 7 2538 247
rect 2542 7 2543 247
rect 2549 7 2550 247
rect 2554 7 2555 247
rect 2561 7 2562 247
rect 2566 7 2567 247
rect 2573 7 2574 247
rect 2578 7 2579 247
rect 2585 7 2586 247
rect 2590 7 2591 247
rect 2597 7 2598 247
rect 2602 7 2603 247
rect 2609 7 2610 247
rect 2614 7 2615 247
rect 2621 7 2622 247
rect 2626 7 2627 247
rect 2633 7 2634 247
rect 2638 7 2639 247
rect 2645 7 2646 247
rect 2650 7 2651 247
rect 2657 7 2658 247
rect 2662 7 2663 247
rect 2669 7 2670 247
rect 2674 7 2675 247
rect 2696 246 2697 250
rect 2694 132 2697 246
rect 2703 244 2709 252
rect 2703 240 2704 244
rect 2708 240 2709 244
rect 2703 132 2709 240
rect 2715 251 2721 252
rect 2715 247 2716 251
rect 2720 247 2721 251
rect 2715 132 2721 247
rect 2727 244 2733 252
rect 2727 240 2728 244
rect 2732 240 2733 244
rect 2727 132 2733 240
rect 2739 245 2742 252
rect 2752 248 2753 252
rect 2739 241 2740 245
rect 2739 132 2742 241
rect 2750 12 2753 248
rect 2759 92 2762 252
rect 2774 245 2777 252
rect 2776 241 2777 245
rect 2774 136 2777 241
rect 2776 132 2777 136
rect 2783 248 2784 252
rect 2796 248 2797 252
rect 2783 136 2786 248
rect 2783 132 2784 136
rect 2794 132 2797 248
rect 2803 132 2809 252
rect 2815 132 2821 252
rect 2827 245 2833 252
rect 2827 241 2828 245
rect 2832 241 2833 245
rect 2827 132 2833 241
rect 2839 250 2842 252
rect 2839 246 2840 250
rect 2839 132 2842 246
rect 2759 88 2760 92
rect 2759 12 2762 88
rect 2859 11 2860 251
rect 2864 11 2865 251
rect 2871 11 2872 251
rect 2876 11 2877 251
rect 2883 11 2884 251
rect 2888 11 2889 251
rect 2895 11 2896 251
rect 2900 11 2901 251
rect 2907 11 2908 251
rect 2912 11 2913 251
rect 2919 11 2920 251
rect 2924 11 2925 251
rect 2931 11 2932 251
rect 2936 11 2937 251
rect 2943 11 2944 251
rect 2948 11 2949 251
rect 2955 11 2956 251
rect 2960 11 2961 251
rect 2967 11 2968 251
rect 2972 11 2973 251
rect 2979 11 2980 251
rect 2984 11 2985 251
rect 2991 11 2992 251
rect 2996 11 2997 251
rect 3003 11 3004 251
rect 3008 11 3009 251
rect 3015 11 3016 251
rect 3020 11 3021 251
rect 3027 11 3028 251
rect 3032 11 3033 251
rect 3039 11 3040 251
rect 3044 11 3045 251
rect 3051 11 3052 251
rect 3056 11 3057 251
rect 3063 11 3064 251
rect 3068 11 3069 251
rect 3075 11 3076 251
rect 3080 11 3081 251
rect 3087 11 3088 251
rect 3092 11 3093 251
rect 3099 11 3100 251
rect 3104 11 3105 251
rect 3111 11 3112 251
rect 3116 11 3117 251
rect 3123 11 3124 251
rect 3128 11 3129 251
rect 3135 11 3136 251
rect 3140 11 3141 251
rect 3147 11 3148 251
rect 3152 11 3153 251
rect 3159 11 3160 251
rect 3164 11 3165 251
rect 3171 11 3172 251
rect 3176 11 3177 251
rect 3183 11 3184 251
rect 3188 11 3189 251
rect 3195 11 3196 251
rect 3200 11 3201 251
rect 3207 11 3208 251
rect 3212 11 3213 251
rect 3219 11 3220 251
rect 3224 11 3225 251
rect 3231 11 3232 251
rect 3236 11 3237 251
rect 3243 11 3244 251
rect 3248 11 3249 251
rect 3255 11 3256 251
rect 3260 11 3261 251
rect 3267 11 3268 251
rect 3272 11 3273 251
rect 3279 11 3280 251
rect 3284 11 3285 251
rect 3291 11 3292 251
rect 3296 11 3297 251
rect 3303 11 3304 251
rect 3308 11 3309 251
rect 3315 11 3316 251
rect 3320 11 3321 251
rect 3327 11 3328 251
rect 3332 11 3333 251
rect 3339 11 3340 251
rect 3344 11 3345 251
rect 3351 11 3352 251
rect 3356 11 3357 251
rect 3363 11 3364 251
rect 3368 11 3369 251
rect 3375 11 3376 251
rect 3380 11 3381 251
rect 3387 11 3388 251
rect 3392 11 3393 251
rect 3399 11 3400 251
rect 3404 11 3405 251
rect 3411 11 3412 251
rect 3416 11 3417 251
rect 3423 11 3424 251
rect 3428 11 3429 251
rect 3435 11 3436 251
rect 3440 11 3441 251
rect 3447 11 3448 251
rect 3452 11 3453 251
rect 3459 11 3460 251
rect 3464 11 3465 251
<< pdiffusion >>
rect 2439 638 2440 642
rect 2442 638 2443 642
rect 2495 638 2496 642
rect 2498 638 2499 642
rect 2428 612 2429 616
rect 2431 612 2432 616
rect 2448 615 2449 619
rect 2451 615 2452 619
rect 2448 607 2449 611
rect 2451 607 2452 611
rect 2549 612 2550 616
rect 2552 612 2556 616
rect 2428 601 2429 605
rect 2431 601 2432 605
rect 2553 610 2556 612
rect 2575 612 2576 616
rect 2578 612 2579 616
rect 2595 612 2596 616
rect 2598 612 2599 616
rect 2560 610 2563 612
rect 2553 606 2557 610
rect 2559 606 2563 610
rect 2553 605 2556 606
rect 2549 601 2550 605
rect 2552 601 2556 605
rect 2428 585 2429 589
rect 2431 585 2432 589
rect 2448 588 2449 592
rect 2451 588 2452 592
rect 2448 580 2449 584
rect 2451 580 2452 584
rect 2549 585 2550 589
rect 2552 585 2556 589
rect 2428 574 2429 578
rect 2431 574 2432 578
rect 2553 583 2556 585
rect 2560 605 2563 606
rect 2575 601 2576 605
rect 2578 601 2579 605
rect 2595 601 2596 605
rect 2598 601 2599 605
rect 2670 610 2674 611
rect 2575 588 2576 592
rect 2578 588 2579 592
rect 2595 588 2596 592
rect 2598 588 2599 592
rect 2560 583 2563 585
rect 2553 579 2557 583
rect 2559 579 2563 583
rect 2670 607 2674 608
rect 2553 578 2556 579
rect 2549 574 2550 578
rect 2552 574 2556 578
rect 2428 558 2429 562
rect 2431 558 2432 562
rect 2448 561 2449 565
rect 2451 561 2452 565
rect 2448 553 2449 557
rect 2451 553 2452 557
rect 2549 558 2550 562
rect 2552 558 2556 562
rect 2428 547 2429 551
rect 2431 547 2432 551
rect 2553 556 2556 558
rect 2560 578 2563 579
rect 2575 577 2576 581
rect 2578 577 2579 581
rect 2595 577 2596 581
rect 2598 577 2599 581
rect 2670 586 2674 587
rect 2575 564 2576 568
rect 2578 564 2579 568
rect 2595 564 2596 568
rect 2598 564 2599 568
rect 2560 556 2563 558
rect 2670 583 2674 584
rect 2553 552 2557 556
rect 2559 552 2563 556
rect 2575 553 2576 557
rect 2578 553 2579 557
rect 2595 553 2596 557
rect 2598 553 2599 557
rect 2553 551 2556 552
rect 2549 547 2550 551
rect 2552 547 2556 551
rect 2428 531 2429 535
rect 2431 531 2432 535
rect 2448 534 2449 538
rect 2451 534 2452 538
rect 2448 526 2449 530
rect 2451 526 2452 530
rect 2549 531 2550 535
rect 2552 531 2556 535
rect 2428 520 2429 524
rect 2431 520 2432 524
rect 2553 529 2556 531
rect 2560 551 2563 552
rect 2670 562 2674 563
rect 2575 540 2576 544
rect 2578 540 2579 544
rect 2595 540 2596 544
rect 2598 540 2599 544
rect 2670 559 2674 560
rect 2560 529 2563 531
rect 2575 529 2576 533
rect 2578 529 2579 533
rect 2595 529 2596 533
rect 2598 529 2599 533
rect 2553 525 2557 529
rect 2559 525 2563 529
rect 2553 524 2556 525
rect 2549 520 2550 524
rect 2552 520 2556 524
rect 2560 524 2563 525
rect 2670 538 2674 539
rect 2670 535 2674 536
rect 2747 533 2750 649
rect 2749 529 2750 533
rect 2756 642 2759 649
rect 2756 638 2757 642
rect 2756 529 2759 638
rect 2820 645 2821 649
rect 2818 529 2821 645
rect 2827 642 2833 649
rect 2827 638 2828 642
rect 2832 638 2833 642
rect 2827 529 2833 638
rect 2839 533 2842 649
rect 2839 529 2840 533
rect 2069 265 2070 505
rect 2074 265 2075 505
rect 2081 265 2082 505
rect 2086 265 2087 505
rect 2093 265 2094 505
rect 2098 265 2099 505
rect 2105 265 2106 505
rect 2110 265 2111 505
rect 2117 265 2118 505
rect 2122 265 2123 505
rect 2129 265 2130 505
rect 2134 265 2135 505
rect 2141 265 2142 505
rect 2146 265 2147 505
rect 2153 265 2154 505
rect 2158 265 2159 505
rect 2165 265 2166 505
rect 2170 265 2171 505
rect 2177 265 2178 505
rect 2182 265 2183 505
rect 2189 265 2190 505
rect 2194 265 2195 505
rect 2201 265 2202 505
rect 2206 265 2207 505
rect 2213 265 2214 505
rect 2218 265 2219 505
rect 2225 265 2226 505
rect 2230 265 2231 505
rect 2237 265 2238 505
rect 2242 265 2243 505
rect 2249 265 2250 505
rect 2254 265 2255 505
rect 2261 265 2262 505
rect 2266 265 2267 505
rect 2273 265 2274 505
rect 2278 265 2279 505
rect 2285 265 2286 505
rect 2290 265 2291 505
rect 2297 265 2298 505
rect 2302 265 2303 505
rect 2309 265 2310 505
rect 2314 265 2315 505
rect 2321 265 2322 505
rect 2326 265 2327 505
rect 2333 265 2334 505
rect 2338 265 2339 505
rect 2345 265 2346 505
rect 2350 265 2351 505
rect 2357 265 2358 505
rect 2362 265 2363 505
rect 2369 265 2370 505
rect 2374 265 2375 505
rect 2381 265 2382 505
rect 2386 265 2387 505
rect 2393 265 2394 505
rect 2398 265 2399 505
rect 2405 265 2406 505
rect 2410 265 2411 505
rect 2417 265 2418 505
rect 2422 265 2423 505
rect 2429 265 2430 505
rect 2434 265 2435 505
rect 2441 265 2442 505
rect 2446 265 2447 505
rect 2453 265 2454 505
rect 2458 265 2459 505
rect 2465 265 2466 505
rect 2470 265 2471 505
rect 2477 265 2478 505
rect 2482 265 2483 505
rect 2489 265 2490 505
rect 2494 265 2495 505
rect 2501 265 2502 505
rect 2506 265 2507 505
rect 2513 265 2514 505
rect 2518 265 2519 505
rect 2525 265 2526 505
rect 2530 265 2531 505
rect 2537 265 2538 505
rect 2542 265 2543 505
rect 2549 265 2550 505
rect 2554 265 2555 505
rect 2561 265 2562 505
rect 2566 265 2567 505
rect 2573 265 2574 505
rect 2578 265 2579 505
rect 2585 265 2586 505
rect 2590 265 2591 505
rect 2597 265 2598 505
rect 2602 265 2603 505
rect 2609 265 2610 505
rect 2614 265 2615 505
rect 2621 265 2622 505
rect 2626 265 2627 505
rect 2633 265 2634 505
rect 2638 265 2639 505
rect 2645 265 2646 505
rect 2650 265 2651 505
rect 2657 265 2658 505
rect 2662 265 2663 505
rect 2669 265 2670 505
rect 2674 265 2675 505
rect 2737 516 2738 520
rect 2735 400 2738 516
rect 2744 516 2745 520
rect 2749 516 2750 520
rect 2744 400 2750 516
rect 2756 411 2759 520
rect 2756 407 2757 411
rect 2756 400 2759 407
rect 2818 404 2821 520
rect 2820 400 2821 404
rect 2827 411 2833 520
rect 2827 407 2828 411
rect 2832 407 2833 411
rect 2827 400 2833 407
rect 2839 516 2840 520
rect 2839 400 2842 516
rect 2696 380 2697 384
rect 2694 270 2697 380
rect 2696 266 2697 270
rect 2694 264 2697 266
rect 2703 275 2709 384
rect 2703 271 2704 275
rect 2708 271 2709 275
rect 2703 264 2709 271
rect 2715 264 2721 384
rect 2727 264 2733 384
rect 2739 268 2742 384
rect 2752 380 2753 384
rect 2750 268 2753 380
rect 2739 264 2740 268
rect 2752 264 2753 268
rect 2759 275 2762 384
rect 2774 275 2777 384
rect 2759 271 2760 275
rect 2776 271 2777 275
rect 2759 264 2762 271
rect 2774 264 2777 271
rect 2783 380 2784 384
rect 2783 268 2786 380
rect 2794 275 2797 384
rect 2796 271 2797 275
rect 2783 264 2784 268
rect 2794 264 2797 271
rect 2803 276 2809 384
rect 2803 272 2804 276
rect 2808 272 2809 276
rect 2803 264 2809 272
rect 2815 269 2821 384
rect 2815 265 2816 269
rect 2820 265 2821 269
rect 2815 264 2821 265
rect 2827 276 2833 384
rect 2827 272 2828 276
rect 2832 272 2833 276
rect 2827 264 2833 272
rect 2839 270 2842 384
rect 2839 266 2840 270
rect 2859 268 2860 508
rect 2864 268 2865 508
rect 2871 268 2872 508
rect 2876 268 2877 508
rect 2883 268 2884 508
rect 2888 268 2889 508
rect 2895 268 2896 508
rect 2900 268 2901 508
rect 2907 268 2908 508
rect 2912 268 2913 508
rect 2919 268 2920 508
rect 2924 268 2925 508
rect 2931 268 2932 508
rect 2936 268 2937 508
rect 2943 268 2944 508
rect 2948 268 2949 508
rect 2955 268 2956 508
rect 2960 268 2961 508
rect 2967 268 2968 508
rect 2972 268 2973 508
rect 2979 268 2980 508
rect 2984 268 2985 508
rect 2991 268 2992 508
rect 2996 268 2997 508
rect 3003 268 3004 508
rect 3008 268 3009 508
rect 3015 268 3016 508
rect 3020 268 3021 508
rect 3027 268 3028 508
rect 3032 268 3033 508
rect 3039 268 3040 508
rect 3044 268 3045 508
rect 3051 268 3052 508
rect 3056 268 3057 508
rect 3063 268 3064 508
rect 3068 268 3069 508
rect 3075 268 3076 508
rect 3080 268 3081 508
rect 3087 268 3088 508
rect 3092 268 3093 508
rect 3099 268 3100 508
rect 3104 268 3105 508
rect 3111 268 3112 508
rect 3116 268 3117 508
rect 3123 268 3124 508
rect 3128 268 3129 508
rect 3135 268 3136 508
rect 3140 268 3141 508
rect 3147 268 3148 508
rect 3152 268 3153 508
rect 3159 268 3160 508
rect 3164 268 3165 508
rect 3171 268 3172 508
rect 3176 268 3177 508
rect 3183 268 3184 508
rect 3188 268 3189 508
rect 3195 268 3196 508
rect 3200 268 3201 508
rect 3207 268 3208 508
rect 3212 268 3213 508
rect 3219 268 3220 508
rect 3224 268 3225 508
rect 3231 268 3232 508
rect 3236 268 3237 508
rect 3243 268 3244 508
rect 3248 268 3249 508
rect 3255 268 3256 508
rect 3260 268 3261 508
rect 3267 268 3268 508
rect 3272 268 3273 508
rect 3279 268 3280 508
rect 3284 268 3285 508
rect 3291 268 3292 508
rect 3296 268 3297 508
rect 3303 268 3304 508
rect 3308 268 3309 508
rect 3315 268 3316 508
rect 3320 268 3321 508
rect 3327 268 3328 508
rect 3332 268 3333 508
rect 3339 268 3340 508
rect 3344 268 3345 508
rect 3351 268 3352 508
rect 3356 268 3357 508
rect 3363 268 3364 508
rect 3368 268 3369 508
rect 3375 268 3376 508
rect 3380 268 3381 508
rect 3387 268 3388 508
rect 3392 268 3393 508
rect 3399 268 3400 508
rect 3404 268 3405 508
rect 3411 268 3412 508
rect 3416 268 3417 508
rect 3423 268 3424 508
rect 3428 268 3429 508
rect 3435 268 3436 508
rect 3440 268 3441 508
rect 3447 268 3448 508
rect 3452 268 3453 508
rect 3459 268 3460 508
rect 3464 268 3465 508
rect 2839 264 2842 266
<< ndcontact >>
rect 2173 687 2177 691
rect 2383 687 2387 691
rect 2796 687 2800 691
rect 2971 687 2975 691
rect 2334 679 2338 683
rect 2544 679 2548 683
rect 2802 679 2806 683
rect 2459 638 2463 642
rect 2467 638 2471 642
rect 2475 638 2479 642
rect 2387 612 2391 616
rect 2402 612 2406 616
rect 2478 615 2482 619
rect 2503 615 2507 619
rect 2387 601 2391 605
rect 2387 585 2391 589
rect 2515 612 2519 616
rect 2523 612 2527 616
rect 2402 601 2406 605
rect 2478 607 2482 611
rect 2503 607 2507 611
rect 2515 601 2519 605
rect 2523 601 2527 605
rect 2402 585 2406 589
rect 2478 588 2482 592
rect 2503 588 2507 592
rect 2387 574 2391 578
rect 2387 558 2391 562
rect 2515 585 2519 589
rect 2523 585 2527 589
rect 2402 574 2406 578
rect 2478 580 2482 584
rect 2503 580 2507 584
rect 2621 612 2625 616
rect 2636 612 2640 616
rect 2654 611 2658 615
rect 2621 601 2625 605
rect 2515 574 2519 578
rect 2523 574 2527 578
rect 2621 588 2625 592
rect 2636 601 2640 605
rect 2654 603 2658 607
rect 2636 588 2640 592
rect 2402 558 2406 562
rect 2478 561 2482 565
rect 2503 561 2507 565
rect 2387 547 2391 551
rect 2387 531 2391 535
rect 2515 558 2519 562
rect 2523 558 2527 562
rect 2402 547 2406 551
rect 2478 553 2482 557
rect 2503 553 2507 557
rect 2654 587 2658 591
rect 2621 577 2625 581
rect 2621 564 2625 568
rect 2636 577 2640 581
rect 2654 579 2658 583
rect 2636 564 2640 568
rect 2515 547 2519 551
rect 2523 547 2527 551
rect 2402 531 2406 535
rect 2478 534 2482 538
rect 2503 534 2507 538
rect 2387 520 2391 524
rect 2515 531 2519 535
rect 2523 531 2527 535
rect 2402 520 2406 524
rect 2478 526 2482 530
rect 2503 526 2507 530
rect 2654 563 2658 567
rect 2621 553 2625 557
rect 2621 540 2625 544
rect 2636 553 2640 557
rect 2654 555 2658 559
rect 2636 540 2640 544
rect 2515 520 2519 524
rect 2523 520 2527 524
rect 2654 539 2658 543
rect 2621 529 2625 533
rect 2636 529 2640 533
rect 2654 531 2658 535
rect 2690 529 2694 533
rect 2702 638 2706 642
rect 2714 645 2718 649
rect 2773 638 2777 642
rect 2785 529 2789 533
rect 2690 516 2694 520
rect 2702 407 2706 411
rect 2714 400 2718 404
rect 2773 407 2777 411
rect 2785 516 2789 520
rect 2797 516 2801 520
rect 2070 7 2074 247
rect 2082 7 2086 247
rect 2094 7 2098 247
rect 2106 7 2110 247
rect 2118 7 2122 247
rect 2130 7 2134 247
rect 2142 7 2146 247
rect 2154 7 2158 247
rect 2166 7 2170 247
rect 2178 7 2182 247
rect 2190 7 2194 247
rect 2202 7 2206 247
rect 2214 7 2218 247
rect 2226 7 2230 247
rect 2238 7 2242 247
rect 2250 7 2254 247
rect 2262 7 2266 247
rect 2274 7 2278 247
rect 2286 7 2290 247
rect 2298 7 2302 247
rect 2310 7 2314 247
rect 2322 7 2326 247
rect 2334 7 2338 247
rect 2346 7 2350 247
rect 2358 7 2362 247
rect 2370 7 2374 247
rect 2382 7 2386 247
rect 2394 7 2398 247
rect 2406 7 2410 247
rect 2418 7 2422 247
rect 2430 7 2434 247
rect 2442 7 2446 247
rect 2454 7 2458 247
rect 2466 7 2470 247
rect 2478 7 2482 247
rect 2490 7 2494 247
rect 2502 7 2506 247
rect 2514 7 2518 247
rect 2526 7 2530 247
rect 2538 7 2542 247
rect 2550 7 2554 247
rect 2562 7 2566 247
rect 2574 7 2578 247
rect 2586 7 2590 247
rect 2598 7 2602 247
rect 2610 7 2614 247
rect 2622 7 2626 247
rect 2634 7 2638 247
rect 2646 7 2650 247
rect 2658 7 2662 247
rect 2670 7 2674 247
rect 2692 246 2696 250
rect 2704 240 2708 244
rect 2716 247 2720 251
rect 2728 240 2732 244
rect 2748 248 2752 252
rect 2740 241 2744 245
rect 2772 241 2776 245
rect 2772 132 2776 136
rect 2784 248 2788 252
rect 2792 248 2796 252
rect 2784 132 2788 136
rect 2828 241 2832 245
rect 2840 246 2844 250
rect 2760 88 2764 92
rect 2860 11 2864 251
rect 2872 11 2876 251
rect 2884 11 2888 251
rect 2896 11 2900 251
rect 2908 11 2912 251
rect 2920 11 2924 251
rect 2932 11 2936 251
rect 2944 11 2948 251
rect 2956 11 2960 251
rect 2968 11 2972 251
rect 2980 11 2984 251
rect 2992 11 2996 251
rect 3004 11 3008 251
rect 3016 11 3020 251
rect 3028 11 3032 251
rect 3040 11 3044 251
rect 3052 11 3056 251
rect 3064 11 3068 251
rect 3076 11 3080 251
rect 3088 11 3092 251
rect 3100 11 3104 251
rect 3112 11 3116 251
rect 3124 11 3128 251
rect 3136 11 3140 251
rect 3148 11 3152 251
rect 3160 11 3164 251
rect 3172 11 3176 251
rect 3184 11 3188 251
rect 3196 11 3200 251
rect 3208 11 3212 251
rect 3220 11 3224 251
rect 3232 11 3236 251
rect 3244 11 3248 251
rect 3256 11 3260 251
rect 3268 11 3272 251
rect 3280 11 3284 251
rect 3292 11 3296 251
rect 3304 11 3308 251
rect 3316 11 3320 251
rect 3328 11 3332 251
rect 3340 11 3344 251
rect 3352 11 3356 251
rect 3364 11 3368 251
rect 3376 11 3380 251
rect 3388 11 3392 251
rect 3400 11 3404 251
rect 3412 11 3416 251
rect 3424 11 3428 251
rect 3436 11 3440 251
rect 3448 11 3452 251
rect 3460 11 3464 251
<< pdcontact >>
rect 2435 638 2439 642
rect 2443 638 2447 642
rect 2491 638 2495 642
rect 2499 638 2503 642
rect 2424 612 2428 616
rect 2432 612 2436 616
rect 2444 615 2448 619
rect 2452 615 2456 619
rect 2444 607 2448 611
rect 2452 607 2456 611
rect 2545 612 2549 616
rect 2424 601 2428 605
rect 2432 601 2436 605
rect 2560 612 2564 616
rect 2571 612 2575 616
rect 2579 612 2583 616
rect 2591 612 2595 616
rect 2599 612 2603 616
rect 2545 601 2549 605
rect 2424 585 2428 589
rect 2432 585 2436 589
rect 2444 588 2448 592
rect 2452 588 2456 592
rect 2444 580 2448 584
rect 2452 580 2456 584
rect 2545 585 2549 589
rect 2424 574 2428 578
rect 2432 574 2436 578
rect 2560 601 2564 605
rect 2571 601 2575 605
rect 2579 601 2583 605
rect 2591 601 2595 605
rect 2599 601 2603 605
rect 2670 611 2674 615
rect 2560 585 2564 589
rect 2571 588 2575 592
rect 2579 588 2583 592
rect 2591 588 2595 592
rect 2599 588 2603 592
rect 2670 603 2674 607
rect 2545 574 2549 578
rect 2424 558 2428 562
rect 2432 558 2436 562
rect 2444 561 2448 565
rect 2452 561 2456 565
rect 2444 553 2448 557
rect 2452 553 2456 557
rect 2545 558 2549 562
rect 2424 547 2428 551
rect 2432 547 2436 551
rect 2560 574 2564 578
rect 2571 577 2575 581
rect 2579 577 2583 581
rect 2591 577 2595 581
rect 2599 577 2603 581
rect 2670 587 2674 591
rect 2571 564 2575 568
rect 2579 564 2583 568
rect 2591 564 2595 568
rect 2599 564 2603 568
rect 2560 558 2564 562
rect 2670 579 2674 583
rect 2571 553 2575 557
rect 2579 553 2583 557
rect 2591 553 2595 557
rect 2599 553 2603 557
rect 2545 547 2549 551
rect 2424 531 2428 535
rect 2432 531 2436 535
rect 2444 534 2448 538
rect 2452 534 2456 538
rect 2444 526 2448 530
rect 2452 526 2456 530
rect 2545 531 2549 535
rect 2424 520 2428 524
rect 2432 520 2436 524
rect 2560 547 2564 551
rect 2670 563 2674 567
rect 2571 540 2575 544
rect 2579 540 2583 544
rect 2591 540 2595 544
rect 2599 540 2603 544
rect 2560 531 2564 535
rect 2670 555 2674 559
rect 2571 529 2575 533
rect 2579 529 2583 533
rect 2591 529 2595 533
rect 2599 529 2603 533
rect 2545 520 2549 524
rect 2670 539 2674 543
rect 2670 531 2674 535
rect 2560 520 2564 524
rect 2745 529 2749 533
rect 2757 638 2761 642
rect 2816 645 2820 649
rect 2828 638 2832 642
rect 2840 529 2844 533
rect 2070 265 2074 505
rect 2082 265 2086 505
rect 2094 265 2098 505
rect 2106 265 2110 505
rect 2118 265 2122 505
rect 2130 265 2134 505
rect 2142 265 2146 505
rect 2154 265 2158 505
rect 2166 265 2170 505
rect 2178 265 2182 505
rect 2190 265 2194 505
rect 2202 265 2206 505
rect 2214 265 2218 505
rect 2226 265 2230 505
rect 2238 265 2242 505
rect 2250 265 2254 505
rect 2262 265 2266 505
rect 2274 265 2278 505
rect 2286 265 2290 505
rect 2298 265 2302 505
rect 2310 265 2314 505
rect 2322 265 2326 505
rect 2334 265 2338 505
rect 2346 265 2350 505
rect 2358 265 2362 505
rect 2370 265 2374 505
rect 2382 265 2386 505
rect 2394 265 2398 505
rect 2406 265 2410 505
rect 2418 265 2422 505
rect 2430 265 2434 505
rect 2442 265 2446 505
rect 2454 265 2458 505
rect 2466 265 2470 505
rect 2478 265 2482 505
rect 2490 265 2494 505
rect 2502 265 2506 505
rect 2514 265 2518 505
rect 2526 265 2530 505
rect 2538 265 2542 505
rect 2550 265 2554 505
rect 2562 265 2566 505
rect 2574 265 2578 505
rect 2586 265 2590 505
rect 2598 265 2602 505
rect 2610 265 2614 505
rect 2622 265 2626 505
rect 2634 265 2638 505
rect 2646 265 2650 505
rect 2658 265 2662 505
rect 2670 265 2674 505
rect 2733 516 2737 520
rect 2745 516 2749 520
rect 2757 407 2761 411
rect 2816 400 2820 404
rect 2828 407 2832 411
rect 2840 516 2844 520
rect 2692 380 2696 384
rect 2692 266 2696 270
rect 2704 271 2708 275
rect 2748 380 2752 384
rect 2740 264 2744 268
rect 2748 264 2752 268
rect 2760 271 2764 275
rect 2772 271 2776 275
rect 2784 380 2788 384
rect 2792 271 2796 275
rect 2784 264 2788 268
rect 2804 272 2808 276
rect 2816 265 2820 269
rect 2828 272 2832 276
rect 2840 266 2844 270
rect 2860 268 2864 508
rect 2872 268 2876 508
rect 2884 268 2888 508
rect 2896 268 2900 508
rect 2908 268 2912 508
rect 2920 268 2924 508
rect 2932 268 2936 508
rect 2944 268 2948 508
rect 2956 268 2960 508
rect 2968 268 2972 508
rect 2980 268 2984 508
rect 2992 268 2996 508
rect 3004 268 3008 508
rect 3016 268 3020 508
rect 3028 268 3032 508
rect 3040 268 3044 508
rect 3052 268 3056 508
rect 3064 268 3068 508
rect 3076 268 3080 508
rect 3088 268 3092 508
rect 3100 268 3104 508
rect 3112 268 3116 508
rect 3124 268 3128 508
rect 3136 268 3140 508
rect 3148 268 3152 508
rect 3160 268 3164 508
rect 3172 268 3176 508
rect 3184 268 3188 508
rect 3196 268 3200 508
rect 3208 268 3212 508
rect 3220 268 3224 508
rect 3232 268 3236 508
rect 3244 268 3248 508
rect 3256 268 3260 508
rect 3268 268 3272 508
rect 3280 268 3284 508
rect 3292 268 3296 508
rect 3304 268 3308 508
rect 3316 268 3320 508
rect 3328 268 3332 508
rect 3340 268 3344 508
rect 3352 268 3356 508
rect 3364 268 3368 508
rect 3376 268 3380 508
rect 3388 268 3392 508
rect 3400 268 3404 508
rect 3412 268 3416 508
rect 3424 268 3428 508
rect 3436 268 3440 508
rect 3448 268 3452 508
rect 3460 268 3464 508
<< psubstratepcontact >>
rect 2395 620 2399 624
rect 2519 620 2523 624
rect 2395 593 2399 597
rect 2519 593 2523 597
rect 2395 566 2399 570
rect 2644 615 2648 619
rect 2644 595 2648 599
rect 2519 566 2523 570
rect 2395 539 2399 543
rect 2644 571 2648 575
rect 2519 539 2523 543
rect 2644 547 2648 551
rect 2684 537 2688 649
rect 2803 524 2807 628
rect 2684 400 2688 512
rect 2803 421 2807 512
rect 2686 130 2690 242
rect 2686 11 2690 126
rect 2766 140 2770 237
rect 2846 129 2850 241
rect 2846 11 2850 125
<< nsubstratencontact >>
rect 2428 620 2432 624
rect 2552 620 2556 624
rect 2428 593 2432 597
rect 2552 593 2556 597
rect 2428 566 2432 570
rect 2670 595 2674 599
rect 2552 566 2556 570
rect 2428 539 2432 543
rect 2670 571 2674 575
rect 2552 539 2556 543
rect 2670 547 2674 551
rect 2727 524 2731 628
rect 2846 537 2850 649
rect 2727 421 2731 512
rect 2846 400 2850 512
rect 2686 274 2690 376
rect 2766 279 2770 387
rect 2846 274 2850 387
<< polysilicon >>
rect 2166 684 2173 686
rect 2338 684 2340 686
rect 2376 684 2383 686
rect 2548 684 2550 686
rect 2789 685 2796 686
rect 2793 684 2796 685
rect 2961 684 2963 686
rect 2968 684 2971 686
rect 3136 685 3142 686
rect 3136 684 3138 685
rect 2695 649 2701 651
rect 2707 649 2713 651
rect 2750 649 2756 651
rect 2778 649 2784 651
rect 2821 649 2827 651
rect 2833 650 2834 651
rect 2838 650 2839 651
rect 2833 649 2839 650
rect 2440 643 2466 645
rect 2440 642 2442 643
rect 2464 642 2466 643
rect 2472 643 2498 645
rect 2472 642 2474 643
rect 2496 642 2498 643
rect 2440 636 2442 638
rect 2392 630 2451 632
rect 2464 633 2466 638
rect 2472 636 2474 638
rect 2496 636 2498 638
rect 2392 611 2394 630
rect 2449 627 2451 630
rect 2477 630 2559 632
rect 2477 627 2479 630
rect 2449 625 2479 627
rect 2449 619 2451 625
rect 2483 619 2491 630
rect 2494 619 2502 622
rect 2399 617 2431 619
rect 2399 616 2401 617
rect 2399 610 2401 612
rect 2409 609 2411 617
rect 2429 616 2431 617
rect 2520 617 2552 619
rect 2520 616 2522 617
rect 2392 584 2394 607
rect 2399 605 2401 607
rect 2429 610 2431 612
rect 2449 611 2451 615
rect 2483 611 2491 615
rect 2494 611 2502 615
rect 2399 600 2401 601
rect 2419 600 2421 608
rect 2520 610 2522 612
rect 2530 609 2532 617
rect 2550 616 2552 617
rect 2429 605 2431 607
rect 2429 600 2431 601
rect 2399 598 2431 600
rect 2449 592 2451 607
rect 2483 592 2491 607
rect 2494 592 2502 607
rect 2520 605 2522 607
rect 2550 610 2552 612
rect 2557 610 2559 630
rect 2576 616 2578 620
rect 2596 617 2628 619
rect 2596 616 2598 617
rect 2520 600 2522 601
rect 2540 600 2542 608
rect 2550 605 2552 607
rect 2550 600 2552 601
rect 2520 598 2552 600
rect 2399 590 2431 592
rect 2399 589 2401 590
rect 2399 583 2401 585
rect 2409 582 2411 590
rect 2429 589 2431 590
rect 2520 590 2552 592
rect 2520 589 2522 590
rect 2392 557 2394 580
rect 2399 578 2401 580
rect 2429 583 2431 585
rect 2449 584 2451 588
rect 2483 584 2491 588
rect 2494 584 2502 588
rect 2399 573 2401 574
rect 2419 573 2421 581
rect 2520 583 2522 585
rect 2530 582 2532 590
rect 2550 589 2552 590
rect 2429 578 2431 580
rect 2429 573 2431 574
rect 2399 571 2431 573
rect 2449 565 2451 580
rect 2483 565 2491 580
rect 2494 565 2502 580
rect 2520 578 2522 580
rect 2550 583 2552 585
rect 2557 583 2559 606
rect 2576 605 2578 612
rect 2596 610 2598 612
rect 2606 609 2608 617
rect 2626 616 2628 617
rect 2596 605 2598 607
rect 2626 610 2628 612
rect 2633 610 2635 634
rect 2576 592 2578 601
rect 2596 600 2598 601
rect 2616 600 2618 608
rect 2626 605 2628 607
rect 2651 608 2654 610
rect 2658 608 2670 610
rect 2674 608 2676 610
rect 2626 600 2628 601
rect 2596 598 2628 600
rect 2596 593 2628 595
rect 2596 592 2598 593
rect 2520 573 2522 574
rect 2540 573 2542 581
rect 2550 578 2552 580
rect 2576 581 2578 588
rect 2596 586 2598 588
rect 2606 585 2608 593
rect 2626 592 2628 593
rect 2596 581 2598 583
rect 2626 586 2628 588
rect 2633 586 2635 606
rect 2550 573 2552 574
rect 2520 571 2552 573
rect 2399 563 2431 565
rect 2399 562 2401 563
rect 2399 556 2401 558
rect 2409 555 2411 563
rect 2429 562 2431 563
rect 2520 563 2552 565
rect 2520 562 2522 563
rect 2392 530 2394 553
rect 2399 551 2401 553
rect 2429 556 2431 558
rect 2449 557 2451 561
rect 2483 557 2491 561
rect 2494 557 2502 561
rect 2399 546 2401 547
rect 2419 546 2421 554
rect 2520 556 2522 558
rect 2530 555 2532 563
rect 2550 562 2552 563
rect 2429 551 2431 553
rect 2429 546 2431 547
rect 2399 544 2431 546
rect 2449 538 2451 553
rect 2483 538 2491 553
rect 2494 538 2502 553
rect 2520 551 2522 553
rect 2550 556 2552 558
rect 2557 556 2559 579
rect 2576 568 2578 577
rect 2596 576 2598 577
rect 2616 576 2618 584
rect 2626 581 2628 583
rect 2651 584 2654 586
rect 2658 584 2670 586
rect 2674 584 2676 586
rect 2626 576 2628 577
rect 2596 574 2628 576
rect 2596 569 2628 571
rect 2596 568 2598 569
rect 2576 557 2578 564
rect 2596 562 2598 564
rect 2606 561 2608 569
rect 2626 568 2628 569
rect 2596 557 2598 559
rect 2626 562 2628 564
rect 2633 562 2635 582
rect 2520 546 2522 547
rect 2540 546 2542 554
rect 2550 551 2552 553
rect 2550 546 2552 547
rect 2520 544 2552 546
rect 2399 536 2431 538
rect 2399 535 2401 536
rect 2399 529 2401 531
rect 2409 528 2411 536
rect 2429 535 2431 536
rect 2520 536 2552 538
rect 2520 535 2522 536
rect 2392 514 2394 526
rect 2399 524 2401 526
rect 2429 529 2431 531
rect 2449 530 2451 534
rect 2483 530 2491 534
rect 2494 530 2502 534
rect 2399 519 2401 520
rect 2419 519 2421 527
rect 2520 529 2522 531
rect 2530 528 2532 536
rect 2550 535 2552 536
rect 2429 524 2431 526
rect 2429 519 2431 520
rect 2399 517 2431 519
rect 2449 514 2451 526
rect 2483 514 2491 526
rect 2494 514 2502 526
rect 2520 524 2522 526
rect 2550 529 2552 531
rect 2557 529 2559 552
rect 2576 544 2578 553
rect 2596 552 2598 553
rect 2616 552 2618 560
rect 2626 557 2628 559
rect 2651 560 2654 562
rect 2658 560 2670 562
rect 2674 560 2676 562
rect 2626 552 2628 553
rect 2596 550 2628 552
rect 2596 545 2628 547
rect 2596 544 2598 545
rect 2576 533 2578 540
rect 2596 538 2598 540
rect 2606 537 2608 545
rect 2626 544 2628 545
rect 2596 533 2598 535
rect 2626 538 2628 540
rect 2633 538 2635 558
rect 2520 519 2522 520
rect 2540 519 2542 527
rect 2550 524 2552 526
rect 2550 519 2552 520
rect 2520 517 2552 519
rect 2557 514 2559 525
rect 2576 524 2578 529
rect 2596 528 2598 529
rect 2616 528 2618 536
rect 2626 533 2628 535
rect 2651 536 2654 538
rect 2658 536 2670 538
rect 2674 536 2676 538
rect 2626 528 2628 529
rect 2596 526 2628 528
rect 2633 524 2635 534
rect 2695 520 2701 529
rect 2707 520 2713 529
rect 2750 528 2756 529
rect 2778 528 2784 529
rect 2750 526 2784 528
rect 2750 522 2784 523
rect 2738 520 2744 522
rect 2750 521 2765 522
rect 2750 520 2756 521
rect 2075 505 2081 508
rect 2087 505 2093 508
rect 2099 505 2105 508
rect 2111 505 2117 508
rect 2123 505 2129 508
rect 2135 505 2141 508
rect 2147 505 2153 508
rect 2159 505 2165 508
rect 2171 505 2177 508
rect 2183 505 2189 508
rect 2195 505 2201 508
rect 2207 505 2213 508
rect 2219 505 2225 508
rect 2231 505 2237 508
rect 2243 505 2249 508
rect 2255 505 2261 508
rect 2267 505 2273 508
rect 2279 505 2285 508
rect 2291 505 2297 508
rect 2303 505 2309 508
rect 2315 505 2321 508
rect 2327 505 2333 508
rect 2339 505 2345 508
rect 2351 505 2357 508
rect 2363 505 2369 508
rect 2375 505 2381 508
rect 2387 505 2393 508
rect 2399 505 2405 508
rect 2411 505 2417 508
rect 2423 505 2429 508
rect 2435 505 2441 508
rect 2447 505 2453 508
rect 2459 505 2465 508
rect 2471 505 2477 508
rect 2483 505 2489 508
rect 2495 505 2501 508
rect 2507 505 2513 508
rect 2519 505 2525 508
rect 2531 505 2537 508
rect 2543 505 2549 508
rect 2555 505 2561 508
rect 2567 505 2573 508
rect 2579 505 2585 508
rect 2591 505 2597 508
rect 2603 505 2609 508
rect 2615 505 2621 508
rect 2627 505 2633 508
rect 2639 505 2645 508
rect 2651 505 2657 508
rect 2663 505 2669 508
rect 1900 262 2066 423
rect 2769 521 2784 522
rect 2778 520 2784 521
rect 2790 520 2796 522
rect 2821 520 2827 529
rect 2833 520 2839 529
rect 2865 508 2871 511
rect 2877 508 2883 511
rect 2889 508 2895 511
rect 2901 508 2907 511
rect 2913 508 2919 511
rect 2925 508 2931 511
rect 2937 508 2943 511
rect 2949 508 2955 511
rect 2961 508 2967 511
rect 2973 508 2979 511
rect 2985 508 2991 511
rect 2997 508 3003 511
rect 3009 508 3015 511
rect 3021 508 3027 511
rect 3033 508 3039 511
rect 3045 508 3051 511
rect 3057 508 3063 511
rect 3069 508 3075 511
rect 3081 508 3087 511
rect 3093 508 3099 511
rect 3105 508 3111 511
rect 3117 508 3123 511
rect 3129 508 3135 511
rect 3141 508 3147 511
rect 3153 508 3159 511
rect 3165 508 3171 511
rect 3177 508 3183 511
rect 3189 508 3195 511
rect 3201 508 3207 511
rect 3213 508 3219 511
rect 3225 508 3231 511
rect 3237 508 3243 511
rect 3249 508 3255 511
rect 3261 508 3267 511
rect 3273 508 3279 511
rect 3285 508 3291 511
rect 3297 508 3303 511
rect 3309 508 3315 511
rect 3321 508 3327 511
rect 3333 508 3339 511
rect 3345 508 3351 511
rect 3357 508 3363 511
rect 3369 508 3375 511
rect 3381 508 3387 511
rect 3393 508 3399 511
rect 3405 508 3411 511
rect 3417 508 3423 511
rect 3429 508 3435 511
rect 3441 508 3447 511
rect 3453 508 3459 511
rect 2695 398 2701 400
rect 2707 399 2713 400
rect 2711 398 2713 399
rect 2738 397 2744 400
rect 2750 398 2756 400
rect 2778 398 2784 400
rect 2790 397 2796 400
rect 2821 399 2827 400
rect 2821 398 2823 399
rect 2833 398 2839 400
rect 2697 385 2734 387
rect 2738 385 2739 387
rect 2697 384 2703 385
rect 2709 384 2715 385
rect 2721 384 2727 385
rect 2733 384 2739 385
rect 2753 384 2759 386
rect 2075 262 2081 265
rect 2087 262 2093 265
rect 2099 262 2105 265
rect 2111 262 2117 265
rect 2123 262 2129 265
rect 2135 262 2141 265
rect 2147 262 2153 265
rect 2159 262 2165 265
rect 2171 262 2177 265
rect 2183 262 2189 265
rect 2195 262 2201 265
rect 2207 262 2213 265
rect 2219 262 2225 265
rect 2231 262 2237 265
rect 2243 262 2249 265
rect 2255 262 2261 265
rect 2267 262 2273 265
rect 2279 262 2285 265
rect 2291 262 2297 265
rect 2303 262 2309 265
rect 2315 262 2321 265
rect 2327 262 2333 265
rect 2339 262 2345 265
rect 2351 262 2357 265
rect 2363 262 2369 265
rect 2375 262 2381 265
rect 2387 262 2393 265
rect 2399 262 2405 265
rect 2411 262 2417 265
rect 2423 262 2429 265
rect 2435 262 2441 265
rect 2447 262 2453 265
rect 2459 262 2465 265
rect 2471 262 2477 265
rect 2483 262 2489 265
rect 2495 262 2501 265
rect 2507 262 2513 265
rect 2519 262 2525 265
rect 2531 262 2537 265
rect 2543 262 2549 265
rect 2555 262 2561 265
rect 2567 262 2573 265
rect 2579 262 2585 265
rect 2591 262 2597 265
rect 2603 262 2609 265
rect 2615 262 2621 265
rect 2627 262 2633 265
rect 2639 262 2645 265
rect 2651 262 2657 265
rect 2663 262 2669 265
rect 2777 384 2783 386
rect 2797 384 2803 386
rect 2809 384 2815 386
rect 2821 384 2827 386
rect 2833 385 2834 386
rect 2838 385 2839 386
rect 2833 384 2839 385
rect 2865 265 2871 268
rect 2877 265 2883 268
rect 2889 265 2895 268
rect 2901 265 2907 268
rect 2913 265 2919 268
rect 2925 265 2931 268
rect 2937 265 2943 268
rect 2949 265 2955 268
rect 2961 265 2967 268
rect 2973 265 2979 268
rect 2985 265 2991 268
rect 2997 265 3003 268
rect 3009 265 3015 268
rect 3021 265 3027 268
rect 3033 265 3039 268
rect 3045 265 3051 268
rect 3057 265 3063 268
rect 3069 265 3075 268
rect 3081 265 3087 268
rect 3093 265 3099 268
rect 3105 265 3111 268
rect 3117 265 3123 268
rect 3129 265 3135 268
rect 3141 265 3147 268
rect 3153 265 3159 268
rect 3165 265 3171 268
rect 3177 265 3183 268
rect 3189 265 3195 268
rect 3201 265 3207 268
rect 3213 265 3219 268
rect 3225 265 3231 268
rect 3237 265 3243 268
rect 3249 265 3255 268
rect 3261 265 3267 268
rect 3273 265 3279 268
rect 3285 265 3291 268
rect 3297 265 3303 268
rect 3309 265 3315 268
rect 3321 265 3327 268
rect 3333 265 3339 268
rect 3345 265 3351 268
rect 3357 265 3363 268
rect 3369 265 3375 268
rect 3381 265 3387 268
rect 3393 265 3399 268
rect 3405 265 3411 268
rect 3417 265 3423 268
rect 3429 265 3435 268
rect 3441 265 3447 268
rect 3453 265 3459 268
rect 3467 265 3633 427
rect 2697 262 2703 264
rect 2709 262 2715 264
rect 2721 262 2727 264
rect 2733 262 2739 264
rect 2753 263 2759 264
rect 2777 263 2783 264
rect 1900 258 2669 262
rect 2753 261 2754 263
rect 2758 261 2783 263
rect 2797 263 2803 264
rect 2809 263 2815 264
rect 2821 263 2827 264
rect 2797 261 2798 263
rect 2802 261 2816 263
rect 2820 261 2827 263
rect 2833 263 2839 264
rect 2833 262 2834 263
rect 2838 262 2839 263
rect 2860 261 3633 265
rect 1900 257 2066 258
rect 2697 253 2698 254
rect 2702 253 2703 254
rect 2697 252 2703 253
rect 2709 253 2716 255
rect 2720 253 2734 255
rect 2738 253 2739 254
rect 2709 252 2715 253
rect 2721 252 2727 253
rect 2733 252 2739 253
rect 2753 253 2778 255
rect 2782 253 2783 255
rect 2753 252 2759 253
rect 2777 252 2783 253
rect 2797 252 2803 254
rect 2809 252 2815 254
rect 2821 252 2827 254
rect 2833 252 2839 254
rect 2075 247 2081 250
rect 2087 247 2093 250
rect 2099 247 2105 250
rect 2111 247 2117 250
rect 2123 247 2129 250
rect 2135 247 2141 250
rect 2147 247 2153 250
rect 2159 247 2165 250
rect 2171 247 2177 250
rect 2183 247 2189 250
rect 2195 247 2201 250
rect 2207 247 2213 250
rect 2219 247 2225 250
rect 2231 247 2237 250
rect 2243 247 2249 250
rect 2255 247 2261 250
rect 2267 247 2273 250
rect 2279 247 2285 250
rect 2291 247 2297 250
rect 2303 247 2309 250
rect 2315 247 2321 250
rect 2327 247 2333 250
rect 2339 247 2345 250
rect 2351 247 2357 250
rect 2363 247 2369 250
rect 2375 247 2381 250
rect 2387 247 2393 250
rect 2399 247 2405 250
rect 2411 247 2417 250
rect 2423 247 2429 250
rect 2435 247 2441 250
rect 2447 247 2453 250
rect 2459 247 2465 250
rect 2471 247 2477 250
rect 2483 247 2489 250
rect 2495 247 2501 250
rect 2507 247 2513 250
rect 2519 247 2525 250
rect 2531 247 2537 250
rect 2543 247 2549 250
rect 2555 247 2561 250
rect 2567 247 2573 250
rect 2579 247 2585 250
rect 2591 247 2597 250
rect 2603 247 2609 250
rect 2615 247 2621 250
rect 2627 247 2633 250
rect 2639 247 2645 250
rect 2651 247 2657 250
rect 2663 247 2669 250
rect 2697 130 2703 132
rect 2709 130 2715 132
rect 2721 130 2727 132
rect 2733 130 2739 132
rect 2865 251 2871 254
rect 2877 251 2883 254
rect 2889 251 2895 254
rect 2901 251 2907 254
rect 2913 251 2919 254
rect 2925 251 2931 254
rect 2937 251 2943 254
rect 2949 251 2955 254
rect 2961 251 2967 254
rect 2973 251 2979 254
rect 2985 251 2991 254
rect 2997 251 3003 254
rect 3009 251 3015 254
rect 3021 251 3027 254
rect 3033 251 3039 254
rect 3045 251 3051 254
rect 3057 251 3063 254
rect 3069 251 3075 254
rect 3081 251 3087 254
rect 3093 251 3099 254
rect 3105 251 3111 254
rect 3117 251 3123 254
rect 3129 251 3135 254
rect 3141 251 3147 254
rect 3153 251 3159 254
rect 3165 251 3171 254
rect 3177 251 3183 254
rect 3189 251 3195 254
rect 3201 251 3207 254
rect 3213 251 3219 254
rect 3225 251 3231 254
rect 3237 251 3243 254
rect 3249 251 3255 254
rect 3261 251 3267 254
rect 3273 251 3279 254
rect 3285 251 3291 254
rect 3297 251 3303 254
rect 3309 251 3315 254
rect 3321 251 3327 254
rect 3333 251 3339 254
rect 3345 251 3351 254
rect 3357 251 3363 254
rect 3369 251 3375 254
rect 3381 251 3387 254
rect 3393 251 3399 254
rect 3405 251 3411 254
rect 3417 251 3423 254
rect 3429 251 3435 254
rect 3441 251 3447 254
rect 3453 251 3459 254
rect 2777 130 2783 132
rect 2797 131 2803 132
rect 2809 131 2815 132
rect 2821 131 2827 132
rect 2833 131 2839 132
rect 2797 129 2798 131
rect 2802 129 2839 131
rect 2753 10 2759 12
rect 2865 8 2871 11
rect 2877 8 2883 11
rect 2889 8 2895 11
rect 2901 8 2907 11
rect 2913 8 2919 11
rect 2925 8 2931 11
rect 2937 8 2943 11
rect 2949 8 2955 11
rect 2961 8 2967 11
rect 2973 8 2979 11
rect 2985 8 2991 11
rect 2997 8 3003 11
rect 3009 8 3015 11
rect 3021 8 3027 11
rect 3033 8 3039 11
rect 3045 8 3051 11
rect 3057 8 3063 11
rect 3069 8 3075 11
rect 3081 8 3087 11
rect 3093 8 3099 11
rect 3105 8 3111 11
rect 3117 8 3123 11
rect 3129 8 3135 11
rect 3141 8 3147 11
rect 3153 8 3159 11
rect 3165 8 3171 11
rect 3177 8 3183 11
rect 3189 8 3195 11
rect 3201 8 3207 11
rect 3213 8 3219 11
rect 3225 8 3231 11
rect 3237 8 3243 11
rect 3249 8 3255 11
rect 3261 8 3267 11
rect 3273 8 3279 11
rect 3285 8 3291 11
rect 3297 8 3303 11
rect 3309 8 3315 11
rect 3321 8 3327 11
rect 3333 8 3339 11
rect 3345 8 3351 11
rect 3357 8 3363 11
rect 3369 8 3375 11
rect 3381 8 3387 11
rect 3393 8 3399 11
rect 3405 8 3411 11
rect 3417 8 3423 11
rect 3429 8 3435 11
rect 3441 8 3447 11
rect 3453 8 3459 11
rect 2075 4 2081 7
rect 2087 4 2093 7
rect 2099 4 2105 7
rect 2111 4 2117 7
rect 2123 4 2129 7
rect 2135 4 2141 7
rect 2147 4 2153 7
rect 2159 4 2165 7
rect 2171 4 2177 7
rect 2183 4 2189 7
rect 2195 4 2201 7
rect 2207 4 2213 7
rect 2219 4 2225 7
rect 2231 4 2237 7
rect 2243 4 2249 7
rect 2255 4 2261 7
rect 2267 4 2273 7
rect 2279 4 2285 7
rect 2291 4 2297 7
rect 2303 4 2309 7
rect 2315 4 2321 7
rect 2327 4 2333 7
rect 2339 4 2345 7
rect 2351 4 2357 7
rect 2363 4 2369 7
rect 2375 4 2381 7
rect 2387 4 2393 7
rect 2399 4 2405 7
rect 2411 4 2417 7
rect 2423 4 2429 7
rect 2435 4 2441 7
rect 2447 4 2453 7
rect 2459 4 2465 7
rect 2471 4 2477 7
rect 2483 4 2489 7
rect 2495 4 2501 7
rect 2507 4 2513 7
rect 2519 4 2525 7
rect 2531 4 2537 7
rect 2543 4 2549 7
rect 2555 4 2561 7
rect 2567 4 2573 7
rect 2579 4 2585 7
rect 2591 4 2597 7
rect 2603 4 2609 7
rect 2615 4 2621 7
rect 2627 4 2633 7
rect 2639 4 2645 7
rect 2651 4 2657 7
rect 2663 4 2669 7
rect 2865 4 3459 8
rect 2075 0 2669 4
<< polycontact >>
rect 2166 680 2170 684
rect 2376 680 2380 684
rect 2789 681 2793 685
rect 3138 681 3142 685
rect 2834 650 2838 654
rect 2451 645 2455 649
rect 2483 645 2487 649
rect 2460 631 2464 635
rect 2631 634 2635 638
rect 2495 622 2499 626
rect 2408 605 2412 609
rect 2418 608 2422 612
rect 2529 605 2533 609
rect 2539 608 2543 612
rect 2575 620 2579 624
rect 2408 578 2412 582
rect 2418 581 2422 585
rect 2529 578 2533 582
rect 2539 581 2543 585
rect 2605 605 2609 609
rect 2615 608 2619 612
rect 2647 608 2651 612
rect 2605 581 2609 585
rect 2615 584 2619 588
rect 2408 551 2412 555
rect 2418 554 2422 558
rect 2529 551 2533 555
rect 2539 554 2543 558
rect 2647 584 2651 588
rect 2605 557 2609 561
rect 2615 560 2619 564
rect 865 518 869 522
rect 2408 524 2412 528
rect 2418 527 2422 531
rect 2529 524 2533 528
rect 2539 527 2543 531
rect 2647 560 2651 564
rect 2605 533 2609 537
rect 2615 536 2619 540
rect 2647 536 2651 540
rect 2765 518 2769 522
rect 2707 395 2711 399
rect 2739 393 2743 397
rect 2791 393 2795 397
rect 2823 395 2827 399
rect 2734 385 2738 389
rect 2834 385 2838 389
rect 2754 259 2758 263
rect 2798 259 2802 263
rect 2816 259 2820 263
rect 2834 259 2838 263
rect 2088 250 2092 254
rect 2100 250 2104 254
rect 2112 250 2116 254
rect 2124 250 2128 254
rect 2136 250 2140 254
rect 2148 250 2152 254
rect 2160 250 2164 254
rect 2172 250 2176 254
rect 2184 250 2188 254
rect 2196 250 2200 254
rect 2208 250 2212 254
rect 2220 250 2224 254
rect 2232 250 2236 254
rect 2244 250 2248 254
rect 2256 250 2260 254
rect 2268 250 2272 254
rect 2280 250 2284 254
rect 2292 250 2296 254
rect 2304 250 2308 254
rect 2316 250 2320 254
rect 2328 250 2332 254
rect 2340 250 2344 254
rect 2352 250 2356 254
rect 2364 250 2368 254
rect 2376 250 2380 254
rect 2388 250 2392 254
rect 2400 250 2404 254
rect 2412 250 2416 254
rect 2424 250 2428 254
rect 2436 250 2440 254
rect 2448 250 2452 254
rect 2460 250 2464 254
rect 2472 250 2476 254
rect 2484 250 2488 254
rect 2496 250 2500 254
rect 2508 250 2512 254
rect 2520 250 2524 254
rect 2532 250 2536 254
rect 2544 250 2548 254
rect 2556 250 2560 254
rect 2568 250 2572 254
rect 2580 250 2584 254
rect 2592 250 2596 254
rect 2604 250 2608 254
rect 2616 250 2620 254
rect 2628 250 2632 254
rect 2640 250 2644 254
rect 2652 250 2656 254
rect 2698 253 2702 257
rect 2716 253 2720 257
rect 2734 253 2738 257
rect 2778 253 2782 257
rect 2798 127 2802 131
<< metal1 >>
rect 2613 708 2814 711
rect 2613 699 2616 708
rect 2723 702 2806 705
rect 2723 699 2726 702
rect 883 691 885 692
rect 865 688 885 691
rect 1933 691 1936 695
rect 2343 691 2346 695
rect 266 654 269 669
rect 865 668 869 688
rect 1933 687 2173 691
rect 2343 687 2383 691
rect 1238 661 1242 669
rect 762 657 1242 661
rect 545 654 593 655
rect 266 652 775 654
rect 266 651 548 652
rect 590 651 771 652
rect 753 618 756 619
rect 735 520 790 524
rect 1686 420 1689 674
rect 1933 667 1936 687
rect 2343 683 2346 687
rect 2166 654 2169 680
rect 2338 680 2346 683
rect 2553 683 2556 695
rect 2613 689 2616 695
rect 2723 688 2726 695
rect 2783 691 2786 695
rect 2765 688 2796 691
rect 2377 664 2380 680
rect 2548 680 2556 683
rect 2765 668 2769 688
rect 2803 683 2806 702
rect 2811 691 2814 708
rect 2811 688 2971 691
rect 2789 677 2792 681
rect 3139 673 3142 681
rect 2789 667 2792 673
rect 3138 661 3142 669
rect 2662 657 3142 661
rect 2445 654 2493 655
rect 2166 652 2675 654
rect 2166 651 2448 652
rect 2490 651 2671 652
rect 2834 649 2838 650
rect 2435 642 2439 645
rect 2467 642 2471 645
rect 2499 642 2503 645
rect 2447 638 2459 642
rect 2479 638 2483 642
rect 2487 638 2491 642
rect 2435 633 2439 638
rect 2392 622 2395 624
rect 2388 620 2395 622
rect 2388 616 2392 620
rect 2432 616 2436 629
rect 2451 625 2455 638
rect 2451 622 2456 625
rect 2453 619 2456 622
rect 2391 612 2392 616
rect 2406 612 2413 616
rect 2417 612 2424 616
rect 2443 615 2444 619
rect 2460 612 2463 631
rect 2467 626 2471 638
rect 2483 626 2487 638
rect 2499 633 2503 638
rect 2483 622 2495 626
rect 2559 624 2563 629
rect 2470 615 2478 619
rect 2507 615 2508 619
rect 2515 616 2519 622
rect 2556 620 2563 624
rect 2575 624 2579 638
rect 2670 631 2677 633
rect 2595 629 2677 631
rect 2591 628 2674 629
rect 2559 616 2563 620
rect 2591 616 2595 628
rect 2639 621 2647 622
rect 2635 619 2647 621
rect 2670 619 2674 628
rect 2635 616 2639 619
rect 2527 612 2534 616
rect 2538 612 2545 616
rect 2559 612 2560 616
rect 2583 612 2584 616
rect 2603 612 2610 616
rect 2614 612 2621 616
rect 2635 612 2636 616
rect 2648 615 2658 619
rect 2388 605 2392 612
rect 2432 605 2436 612
rect 2452 611 2463 612
rect 2443 607 2444 611
rect 2456 609 2463 611
rect 2470 608 2478 611
rect 2507 607 2508 611
rect 2391 601 2392 605
rect 2406 601 2413 605
rect 2417 601 2424 605
rect 2388 597 2392 601
rect 2388 593 2395 597
rect 2388 589 2392 593
rect 2432 589 2436 601
rect 2453 602 2459 604
rect 2515 605 2519 612
rect 2559 605 2563 612
rect 2591 605 2595 612
rect 2635 605 2639 612
rect 2670 615 2681 619
rect 2453 601 2462 602
rect 2466 601 2502 604
rect 2453 592 2456 601
rect 2466 598 2469 601
rect 2527 601 2534 605
rect 2538 601 2545 605
rect 2559 601 2560 605
rect 2583 601 2584 605
rect 2603 601 2610 605
rect 2614 601 2621 605
rect 2635 601 2636 605
rect 2658 603 2666 607
rect 2391 585 2392 589
rect 2406 585 2413 589
rect 2417 585 2424 589
rect 2443 588 2444 592
rect 2460 595 2469 598
rect 2460 585 2463 595
rect 2470 588 2478 592
rect 2507 588 2508 592
rect 2515 589 2519 601
rect 2559 597 2563 601
rect 2556 593 2563 597
rect 2559 589 2563 593
rect 2591 592 2595 601
rect 2635 598 2639 601
rect 2677 599 2681 615
rect 2635 595 2644 598
rect 2648 595 2658 599
rect 2674 595 2681 599
rect 2635 592 2639 595
rect 2527 585 2534 589
rect 2538 585 2545 589
rect 2559 585 2560 589
rect 2583 588 2584 592
rect 2603 588 2610 592
rect 2614 588 2621 592
rect 2635 588 2636 592
rect 2654 591 2658 595
rect 2677 591 2681 595
rect 2388 578 2392 585
rect 2432 578 2436 585
rect 2452 584 2463 585
rect 2443 580 2444 584
rect 2456 582 2463 584
rect 2470 581 2478 584
rect 2507 580 2508 584
rect 2391 574 2392 578
rect 2406 574 2413 578
rect 2417 574 2424 578
rect 2388 570 2392 574
rect 2388 566 2395 570
rect 2388 562 2392 566
rect 2432 562 2436 574
rect 2453 575 2459 577
rect 2515 578 2519 585
rect 2559 578 2563 585
rect 2591 581 2595 588
rect 2635 581 2639 588
rect 2674 587 2681 591
rect 2453 574 2462 575
rect 2466 574 2502 577
rect 2453 565 2456 574
rect 2466 571 2469 574
rect 2527 574 2534 578
rect 2538 574 2545 578
rect 2559 574 2560 578
rect 2583 577 2584 581
rect 2603 577 2610 581
rect 2614 577 2621 581
rect 2635 577 2636 581
rect 2658 579 2666 583
rect 2391 558 2392 562
rect 2406 558 2413 562
rect 2417 558 2424 562
rect 2443 561 2444 565
rect 2460 568 2469 571
rect 2460 558 2463 568
rect 2470 561 2478 565
rect 2507 561 2508 565
rect 2515 562 2519 574
rect 2559 570 2563 574
rect 2556 566 2563 570
rect 2591 568 2595 577
rect 2635 574 2639 577
rect 2677 575 2681 587
rect 2635 571 2644 574
rect 2648 571 2658 575
rect 2674 571 2681 575
rect 2635 568 2639 571
rect 2559 562 2563 566
rect 2583 564 2584 568
rect 2603 564 2610 568
rect 2614 564 2621 568
rect 2635 564 2636 568
rect 2654 567 2658 571
rect 2677 567 2681 571
rect 2527 558 2534 562
rect 2538 558 2545 562
rect 2559 558 2560 562
rect 2388 551 2392 558
rect 2432 551 2436 558
rect 2452 557 2463 558
rect 2443 553 2444 557
rect 2456 555 2463 557
rect 2470 554 2478 557
rect 2507 553 2508 557
rect 2391 547 2392 551
rect 2406 547 2413 551
rect 2417 547 2424 551
rect 2388 543 2392 547
rect 2388 539 2395 543
rect 2388 535 2392 539
rect 2432 535 2436 547
rect 2453 548 2459 550
rect 2515 551 2519 558
rect 2559 551 2563 558
rect 2591 557 2595 564
rect 2635 557 2639 564
rect 2674 563 2681 567
rect 2583 553 2584 557
rect 2603 553 2610 557
rect 2614 553 2621 557
rect 2635 553 2636 557
rect 2658 555 2666 559
rect 2453 547 2462 548
rect 2466 547 2502 550
rect 2453 538 2456 547
rect 2466 544 2469 547
rect 2527 547 2534 551
rect 2538 547 2545 551
rect 2559 547 2560 551
rect 2391 531 2392 535
rect 2406 531 2413 535
rect 2417 531 2424 535
rect 2443 534 2444 538
rect 2460 541 2469 544
rect 2460 531 2463 541
rect 2470 534 2478 538
rect 2507 534 2508 538
rect 2515 535 2519 547
rect 2559 543 2563 547
rect 2591 544 2595 553
rect 2635 550 2639 553
rect 2677 551 2681 563
rect 2635 547 2644 550
rect 2648 547 2658 551
rect 2674 547 2681 551
rect 2635 544 2639 547
rect 2556 539 2563 543
rect 2583 540 2584 544
rect 2603 540 2610 544
rect 2614 540 2621 544
rect 2635 540 2636 544
rect 2654 543 2658 547
rect 2677 543 2681 547
rect 2559 535 2563 539
rect 2527 531 2534 535
rect 2538 531 2545 535
rect 2559 531 2560 535
rect 2591 533 2595 540
rect 2635 533 2639 540
rect 2674 539 2681 543
rect 2718 645 2816 649
rect 2820 645 2838 649
rect 2706 638 2757 642
rect 2777 638 2828 642
rect 2727 631 2846 635
rect 2727 628 2731 631
rect 2388 524 2392 531
rect 2432 524 2436 531
rect 2452 530 2463 531
rect 2443 526 2444 530
rect 2456 528 2463 530
rect 2470 527 2478 530
rect 2507 526 2508 530
rect 2391 520 2392 524
rect 2406 520 2413 524
rect 2417 520 2424 524
rect 2388 514 2392 520
rect 2432 514 2436 520
rect 2453 521 2459 523
rect 2515 524 2519 531
rect 2559 524 2563 531
rect 2583 529 2584 533
rect 2603 529 2610 533
rect 2614 529 2621 533
rect 2635 529 2636 533
rect 2658 531 2666 535
rect 2684 533 2688 537
rect 2684 529 2690 533
rect 2591 524 2595 529
rect 2635 524 2639 529
rect 2690 524 2694 529
rect 2453 520 2462 521
rect 2466 520 2502 523
rect 2453 514 2456 520
rect 2466 517 2469 520
rect 2527 520 2534 524
rect 2538 520 2545 524
rect 2559 520 2560 524
rect 2635 520 2694 524
rect 2460 514 2469 517
rect 2515 514 2519 520
rect 2559 514 2563 520
rect 2684 516 2690 520
rect 2727 520 2731 524
rect 2745 520 2749 529
rect 2727 516 2733 520
rect 2785 520 2789 529
rect 2846 533 2850 537
rect 2803 520 2807 524
rect 2801 516 2807 520
rect 2844 529 2850 533
rect 2840 520 2844 529
rect 2844 516 2850 520
rect 2684 512 2688 516
rect 2082 508 2662 511
rect 2082 505 2086 508
rect 2106 505 2110 508
rect 2130 505 2134 508
rect 2154 505 2158 508
rect 2178 505 2182 508
rect 2202 505 2206 508
rect 2226 505 2230 508
rect 2250 505 2254 508
rect 2274 505 2278 508
rect 2298 505 2302 508
rect 2322 505 2326 508
rect 2346 505 2350 508
rect 2370 505 2374 508
rect 2394 505 2398 508
rect 2418 505 2422 508
rect 2442 505 2446 508
rect 2466 505 2470 508
rect 2490 505 2494 508
rect 2514 505 2518 508
rect 2538 505 2542 508
rect 2562 505 2566 508
rect 2586 505 2590 508
rect 2610 505 2614 508
rect 2634 505 2638 508
rect 2658 505 2662 508
rect 2055 262 2059 264
rect 2727 512 2731 516
rect 2803 512 2807 516
rect 2803 418 2807 421
rect 2688 414 2807 418
rect 2846 515 2850 516
rect 2846 512 3452 515
rect 2706 407 2757 411
rect 2777 407 2828 411
rect 2718 400 2816 404
rect 2850 511 3452 512
rect 2872 508 2876 511
rect 2896 508 2900 511
rect 2920 508 2924 511
rect 2944 508 2948 511
rect 2968 508 2972 511
rect 2992 508 2996 511
rect 3016 508 3020 511
rect 3040 508 3044 511
rect 3064 508 3068 511
rect 3088 508 3092 511
rect 3112 508 3116 511
rect 3136 508 3140 511
rect 3160 508 3164 511
rect 3184 508 3188 511
rect 3208 508 3212 511
rect 3232 508 3236 511
rect 3256 508 3260 511
rect 3280 508 3284 511
rect 3304 508 3308 511
rect 3328 508 3332 511
rect 3352 508 3356 511
rect 3376 508 3380 511
rect 3400 508 3404 511
rect 3424 508 3428 511
rect 3448 508 3452 511
rect 2707 393 2711 395
rect 2692 389 2711 393
rect 2739 389 2743 393
rect 2784 389 2795 393
rect 2823 394 2827 395
rect 2823 390 2838 394
rect 2834 389 2838 390
rect 2692 384 2696 389
rect 2738 385 2752 389
rect 2748 384 2752 385
rect 2674 372 2686 376
rect 2690 279 2708 283
rect 2704 275 2708 279
rect 2784 384 2788 389
rect 2766 275 2770 279
rect 2792 279 2846 283
rect 2792 275 2796 279
rect 2708 271 2760 275
rect 2764 271 2772 275
rect 2776 271 2792 275
rect 2808 272 2828 276
rect 2070 262 2074 265
rect 2094 262 2098 265
rect 2118 262 2122 265
rect 2142 262 2146 265
rect 2166 262 2170 265
rect 2190 262 2194 265
rect 2214 262 2218 265
rect 2238 262 2242 265
rect 2262 262 2266 265
rect 2286 262 2290 265
rect 2310 262 2314 265
rect 2334 262 2338 265
rect 2358 262 2362 265
rect 2382 262 2386 265
rect 2406 262 2410 265
rect 2430 262 2434 265
rect 2454 262 2458 265
rect 2478 262 2482 265
rect 2502 262 2506 265
rect 2526 262 2530 265
rect 2550 262 2554 265
rect 2574 262 2578 265
rect 2598 262 2602 265
rect 2622 262 2626 265
rect 2646 262 2650 265
rect 2670 262 2674 265
rect 2055 258 2674 262
rect 2082 254 2662 258
rect 2082 250 2088 254
rect 2092 250 2100 254
rect 2104 250 2112 254
rect 2116 250 2124 254
rect 2128 250 2136 254
rect 2140 250 2148 254
rect 2152 250 2160 254
rect 2164 250 2172 254
rect 2176 250 2184 254
rect 2188 250 2196 254
rect 2200 250 2208 254
rect 2212 250 2220 254
rect 2224 250 2232 254
rect 2236 250 2244 254
rect 2248 250 2256 254
rect 2260 250 2268 254
rect 2272 250 2280 254
rect 2284 250 2292 254
rect 2296 250 2304 254
rect 2308 250 2316 254
rect 2320 250 2328 254
rect 2332 250 2340 254
rect 2344 250 2352 254
rect 2356 250 2364 254
rect 2368 250 2376 254
rect 2380 250 2388 254
rect 2392 250 2400 254
rect 2404 250 2412 254
rect 2416 250 2424 254
rect 2428 250 2436 254
rect 2440 250 2448 254
rect 2452 250 2460 254
rect 2464 250 2472 254
rect 2476 250 2484 254
rect 2488 250 2496 254
rect 2500 250 2508 254
rect 2512 250 2520 254
rect 2524 250 2532 254
rect 2536 250 2544 254
rect 2548 250 2556 254
rect 2560 250 2568 254
rect 2572 250 2580 254
rect 2584 250 2592 254
rect 2596 250 2604 254
rect 2608 250 2616 254
rect 2620 250 2628 254
rect 2632 250 2640 254
rect 2644 250 2652 254
rect 2656 250 2662 254
rect 2082 247 2086 250
rect 2106 247 2110 250
rect 2130 247 2134 250
rect 2154 247 2158 250
rect 2178 247 2182 250
rect 2202 247 2206 250
rect 2226 247 2230 250
rect 2250 247 2254 250
rect 2274 247 2278 250
rect 2298 247 2302 250
rect 2322 247 2326 250
rect 2346 247 2350 250
rect 2370 247 2374 250
rect 2394 247 2398 250
rect 2418 247 2422 250
rect 2442 247 2446 250
rect 2466 247 2470 250
rect 2490 247 2494 250
rect 2514 247 2518 250
rect 2538 247 2542 250
rect 2562 247 2566 250
rect 2586 247 2590 250
rect 2610 247 2614 250
rect 2634 247 2638 250
rect 2658 247 2662 250
rect 2692 257 2696 266
rect 2740 257 2744 264
rect 2692 253 2698 257
rect 2738 253 2744 257
rect 2748 263 2752 264
rect 2748 259 2754 263
rect 2692 250 2696 253
rect 2716 251 2720 253
rect 2748 252 2752 259
rect 2784 257 2788 264
rect 2816 263 2820 265
rect 2840 263 2844 266
rect 2782 253 2788 257
rect 2784 252 2788 253
rect 2792 259 2798 263
rect 2838 259 2844 263
rect 3586 420 3589 695
rect 2860 265 2864 268
rect 2884 265 2888 268
rect 2908 265 2912 268
rect 2932 265 2936 268
rect 2956 265 2960 268
rect 2980 265 2984 268
rect 3004 265 3008 268
rect 3028 265 3032 268
rect 3052 265 3056 268
rect 3076 265 3080 268
rect 3100 265 3104 268
rect 3124 265 3128 268
rect 3148 265 3152 268
rect 3172 265 3176 268
rect 3196 265 3200 268
rect 3220 265 3224 268
rect 3244 265 3248 268
rect 3268 265 3272 268
rect 3292 265 3296 268
rect 3316 265 3320 268
rect 3340 265 3344 268
rect 3364 265 3368 268
rect 3388 265 3392 268
rect 3412 265 3416 268
rect 3436 265 3440 268
rect 3460 265 3464 268
rect 3474 265 3478 270
rect 2860 261 3478 265
rect 2792 252 2796 259
rect 2840 250 2844 259
rect 2865 258 3459 261
rect 2872 254 3452 258
rect 2872 251 2876 254
rect 2896 251 2900 254
rect 2920 251 2924 254
rect 2944 251 2948 254
rect 2968 251 2972 254
rect 2992 251 2996 254
rect 3016 251 3020 254
rect 3040 251 3044 254
rect 3064 251 3068 254
rect 3088 251 3092 254
rect 3112 251 3116 254
rect 3136 251 3140 254
rect 3160 251 3164 254
rect 3184 251 3188 254
rect 3208 251 3212 254
rect 3232 251 3236 254
rect 3256 251 3260 254
rect 3280 251 3284 254
rect 3304 251 3308 254
rect 3328 251 3332 254
rect 3352 251 3356 254
rect 3376 251 3380 254
rect 3400 251 3404 254
rect 3424 251 3428 254
rect 3448 251 3452 254
rect 2070 4 2074 7
rect 2094 4 2098 7
rect 2118 4 2122 7
rect 2142 4 2146 7
rect 2166 4 2170 7
rect 2190 4 2194 7
rect 2214 4 2218 7
rect 2238 4 2242 7
rect 2262 4 2266 7
rect 2286 4 2290 7
rect 2310 4 2314 7
rect 2334 4 2338 7
rect 2358 4 2362 7
rect 2382 4 2386 7
rect 2406 4 2410 7
rect 2430 4 2434 7
rect 2454 4 2458 7
rect 2478 4 2482 7
rect 2502 4 2506 7
rect 2526 4 2530 7
rect 2550 4 2554 7
rect 2574 4 2578 7
rect 2598 4 2602 7
rect 2622 4 2626 7
rect 2646 4 2650 7
rect 2670 4 2674 7
rect 2708 240 2728 244
rect 2744 241 2772 245
rect 2776 241 2828 245
rect 2740 237 2744 241
rect 2690 233 2744 237
rect 2766 237 2770 241
rect 2828 237 2832 241
rect 2828 233 2846 237
rect 2766 136 2770 140
rect 2766 132 2772 136
rect 2686 126 2690 130
rect 2772 124 2776 132
rect 2784 131 2788 132
rect 2784 127 2798 131
rect 2846 125 2850 129
rect 2772 120 2773 124
rect 2764 88 2773 92
rect 2686 4 2690 11
rect 2846 8 2850 11
rect 2860 8 2864 11
rect 2884 8 2888 11
rect 2908 8 2912 11
rect 2932 8 2936 11
rect 2956 8 2960 11
rect 2980 8 2984 11
rect 3004 8 3008 11
rect 3028 8 3032 11
rect 3052 8 3056 11
rect 3076 8 3080 11
rect 3100 8 3104 11
rect 3124 8 3128 11
rect 3148 8 3152 11
rect 3172 8 3176 11
rect 3196 8 3200 11
rect 3220 8 3224 11
rect 3244 8 3248 11
rect 3268 8 3272 11
rect 3292 8 3296 11
rect 3316 8 3320 11
rect 3340 8 3344 11
rect 3364 8 3368 11
rect 3388 8 3392 11
rect 3412 8 3416 11
rect 3436 8 3440 11
rect 3460 8 3464 11
rect 2846 4 3464 8
rect 2070 0 2690 4
<< m2contact >>
rect 889 673 893 677
rect 480 664 484 668
rect 865 664 869 668
rect 1238 669 1242 673
rect 758 657 762 661
rect 771 648 775 652
rect 823 625 827 629
rect 766 603 770 607
rect 766 579 770 583
rect 766 555 770 559
rect 766 531 770 535
rect 865 522 869 526
rect 2380 664 2384 668
rect 2765 664 2769 668
rect 2789 673 2793 677
rect 3138 669 3142 673
rect 2658 657 2662 661
rect 2671 648 2675 652
rect 2483 638 2487 642
rect 2432 629 2439 633
rect 2388 622 2392 626
rect 2413 612 2417 616
rect 2439 615 2443 619
rect 2467 622 2471 626
rect 2575 638 2579 642
rect 2499 629 2503 633
rect 2559 629 2563 633
rect 2515 622 2519 626
rect 2466 615 2470 619
rect 2508 615 2512 619
rect 2631 638 2635 642
rect 2591 629 2595 633
rect 2677 629 2681 633
rect 2635 621 2639 625
rect 2534 612 2538 616
rect 2567 612 2571 616
rect 2584 612 2588 616
rect 2610 612 2614 616
rect 2439 607 2443 611
rect 2466 608 2470 612
rect 2508 607 2512 611
rect 2413 601 2417 605
rect 2459 602 2463 606
rect 2643 608 2647 612
rect 2502 600 2506 604
rect 2534 601 2538 605
rect 2567 601 2571 605
rect 2584 601 2588 605
rect 2610 601 2614 605
rect 2666 603 2670 607
rect 2413 585 2417 589
rect 2439 588 2443 592
rect 2466 588 2470 592
rect 2508 588 2512 592
rect 2534 585 2538 589
rect 2567 588 2571 592
rect 2584 588 2588 592
rect 2610 588 2614 592
rect 2439 580 2443 584
rect 2466 581 2470 585
rect 2508 580 2512 584
rect 2413 574 2417 578
rect 2459 575 2463 579
rect 2643 584 2647 588
rect 2502 573 2506 577
rect 2534 574 2538 578
rect 2567 577 2571 581
rect 2584 577 2588 581
rect 2610 577 2614 581
rect 2666 579 2670 583
rect 2413 558 2417 562
rect 2439 561 2443 565
rect 2466 561 2470 565
rect 2508 561 2512 565
rect 2567 564 2571 568
rect 2584 564 2588 568
rect 2610 564 2614 568
rect 2534 558 2538 562
rect 2439 553 2443 557
rect 2466 554 2470 558
rect 2508 553 2512 557
rect 2413 547 2417 551
rect 2459 548 2463 552
rect 2643 560 2647 564
rect 2567 553 2571 557
rect 2584 553 2588 557
rect 2610 553 2614 557
rect 2666 555 2670 559
rect 2502 546 2506 550
rect 2534 547 2538 551
rect 2413 531 2417 535
rect 2439 534 2443 538
rect 2466 534 2470 538
rect 2508 534 2512 538
rect 2567 540 2571 544
rect 2584 540 2588 544
rect 2610 540 2614 544
rect 2534 531 2538 535
rect 2643 536 2647 540
rect 2723 625 2727 629
rect 2439 526 2443 530
rect 2466 527 2470 531
rect 2508 526 2512 530
rect 2413 520 2417 524
rect 2459 521 2463 525
rect 2567 529 2571 533
rect 2584 529 2588 533
rect 2610 529 2614 533
rect 2666 531 2670 535
rect 2502 519 2506 523
rect 2534 520 2538 524
rect 2765 522 2769 526
<< metal2 >>
rect 765 673 889 674
rect 2665 673 2789 674
rect 765 671 892 673
rect 484 664 749 667
rect 746 636 749 664
rect 746 633 756 636
rect 753 607 756 633
rect 759 614 762 657
rect 765 620 768 671
rect 2665 671 2792 673
rect 2384 664 2649 667
rect 771 626 774 648
rect 777 629 786 633
rect 771 623 776 626
rect 782 625 823 629
rect 765 617 770 620
rect 759 611 763 614
rect 752 604 756 607
rect 752 576 755 604
rect 760 600 763 611
rect 767 607 770 617
rect 760 597 769 600
rect 766 583 769 597
rect 752 573 769 576
rect 766 559 769 573
rect 773 535 776 623
rect 770 532 776 535
rect 865 526 869 664
rect 2487 639 2575 642
rect 2579 639 2631 642
rect 2646 636 2649 664
rect 2646 633 2656 636
rect 2439 629 2499 633
rect 2503 629 2559 633
rect 2563 629 2591 633
rect 2392 622 2467 626
rect 2471 622 2515 626
rect 2519 622 2635 626
rect 2413 616 2439 619
rect 2443 616 2466 619
rect 2493 615 2508 618
rect 2512 616 2522 619
rect 2512 615 2534 616
rect 2420 611 2466 612
rect 2420 609 2439 611
rect 2420 605 2423 609
rect 2443 609 2466 611
rect 2417 601 2423 605
rect 2493 605 2496 615
rect 2519 612 2534 615
rect 2538 612 2567 616
rect 2588 612 2610 616
rect 2463 602 2496 605
rect 2512 605 2515 611
rect 2610 608 2643 612
rect 2653 607 2656 633
rect 2659 614 2662 657
rect 2665 620 2668 671
rect 2671 626 2674 648
rect 2681 629 2686 633
rect 2671 623 2676 626
rect 2682 625 2723 629
rect 2665 617 2670 620
rect 2659 611 2663 614
rect 2512 604 2534 605
rect 2506 601 2534 604
rect 2538 601 2567 605
rect 2588 601 2610 605
rect 2652 604 2656 607
rect 2413 589 2439 592
rect 2443 589 2466 592
rect 2493 588 2508 591
rect 2512 589 2522 592
rect 2534 589 2567 592
rect 2512 588 2534 589
rect 2420 584 2466 585
rect 2420 582 2439 584
rect 2420 578 2423 582
rect 2443 582 2466 584
rect 2417 574 2423 578
rect 2493 578 2496 588
rect 2519 585 2534 588
rect 2538 588 2567 589
rect 2588 588 2610 592
rect 2610 584 2643 588
rect 2463 575 2496 578
rect 2512 578 2515 584
rect 2534 578 2567 581
rect 2512 577 2534 578
rect 2506 574 2534 577
rect 2538 577 2567 578
rect 2588 577 2610 581
rect 2652 576 2655 604
rect 2660 600 2663 611
rect 2667 607 2670 617
rect 2660 597 2669 600
rect 2666 583 2669 597
rect 2652 573 2669 576
rect 2413 562 2439 565
rect 2443 562 2466 565
rect 2493 561 2508 564
rect 2512 562 2522 565
rect 2534 564 2567 568
rect 2588 564 2610 568
rect 2534 562 2538 564
rect 2512 561 2534 562
rect 2420 557 2466 558
rect 2420 555 2439 557
rect 2420 551 2423 555
rect 2443 555 2466 557
rect 2417 547 2423 551
rect 2493 551 2496 561
rect 2519 558 2534 561
rect 2610 560 2643 564
rect 2666 559 2669 573
rect 2463 548 2496 551
rect 2512 551 2515 557
rect 2588 553 2610 557
rect 2567 551 2571 553
rect 2512 550 2534 551
rect 2506 547 2534 550
rect 2538 547 2571 551
rect 2534 540 2567 544
rect 2588 540 2610 544
rect 2413 535 2439 538
rect 2443 535 2466 538
rect 2493 534 2508 537
rect 2512 535 2522 538
rect 2534 535 2538 540
rect 2610 536 2643 540
rect 2673 535 2676 623
rect 2512 534 2534 535
rect 2420 530 2466 531
rect 2420 528 2439 530
rect 2420 524 2423 528
rect 2443 528 2466 530
rect 2417 520 2423 524
rect 2493 524 2496 534
rect 2519 531 2534 534
rect 2463 521 2496 524
rect 2512 524 2515 530
rect 2588 529 2610 533
rect 2670 532 2676 535
rect 2567 524 2571 529
rect 2512 523 2534 524
rect 2506 520 2534 523
rect 2538 520 2571 524
rect 2765 526 2769 664
<< high_resist >>
rect 1940 700 2340 702
rect 2350 700 2550 702
rect 2560 700 2610 702
rect 2620 700 2720 702
rect 2730 700 2780 702
rect 2791 700 3583 702
rect 1940 693 2340 695
rect 2350 693 2550 695
rect 2560 693 2610 695
rect 2620 693 2720 695
rect 2730 693 2780 695
rect 2791 693 3583 695
rect 2770 94 2772 118
rect 2778 94 2780 118
<< poly2_high_resist >>
rect 1940 695 2340 700
rect 2350 695 2550 700
rect 2560 695 2610 700
rect 2620 695 2720 700
rect 2730 695 2780 700
rect 2791 695 3583 700
rect 2772 94 2778 118
use resistors  resistors_0
timestamp 1418855221
transform -1 0 1688 0 -1 699
box -3 -12 1656 35
use spi-interface  spi-interface_0
timestamp 1418856619
transform 0 1 502 -1 0 622
box -27 -21 108 279
use amplifier  amplifier_0
timestamp 1418853988
transform 1 0 781 0 1 394
box -781 -394 952 261
use chip  chip_0
timestamp 1259953556
transform 1 0 -709 0 1 -751
box 0 0 5000 5000
<< labels >>
rlabel metal2 765 634 768 636 1 B0
rlabel metal2 759 634 762 636 1 B1
rlabel metal2 753 634 756 636 1 B2
rlabel metal2 771 634 774 636 1 B3
rlabel metal2 2665 634 2668 636 1 B0
rlabel metal2 2659 634 2662 636 1 B1
rlabel metal2 2653 634 2656 636 1 B2
rlabel metal2 2671 634 2674 636 1 B3
rlabel metal1 2789 667 2792 675 5 B0
rlabel metal1 2377 664 2380 674 1 B2
rlabel metal1 2166 669 2169 680 5 B3
rlabel metal1 1933 667 1936 695 3 Vref
rlabel metal1 3139 673 3142 681 5 B1
rlabel metal1 3586 667 3589 695 7 Vout
rlabel metal2 2402 622 2406 626 3 Gnd
rlabel m2contact 2591 629 2595 633 3 Vdd
rlabel metal1 2635 547 2639 548 6 Gnd
rlabel metal1 2591 524 2595 525 1 Vdd
rlabel m2contact 2584 540 2588 544 7 Qbar
rlabel pdcontact 2571 540 2575 544 7 Dbar
rlabel m2contact 2584 529 2588 533 1 Q
rlabel pdcontact 2571 529 2575 533 1 D
rlabel polysilicon 2576 524 2578 525 1 En
rlabel polysilicon 2633 524 2635 525 1 En
rlabel metal1 2662 531 2666 535 7 Qout
rlabel pdcontact 2670 539 2674 543 7 Vdd
rlabel ndcontact 2654 539 2658 543 3 Gnd
rlabel metal1 2635 571 2639 572 6 Gnd
rlabel metal1 2591 548 2595 549 1 Vdd
rlabel m2contact 2584 564 2588 568 7 Qbar
rlabel pdcontact 2571 564 2575 568 7 Dbar
rlabel m2contact 2584 553 2588 557 1 Q
rlabel pdcontact 2571 553 2575 557 1 D
rlabel polysilicon 2576 548 2578 549 1 En
rlabel polysilicon 2633 548 2635 549 1 En
rlabel metal1 2662 555 2666 559 7 Qout
rlabel pdcontact 2670 563 2674 567 7 Vdd
rlabel ndcontact 2654 563 2658 567 3 Gnd
rlabel metal1 2635 595 2639 596 6 Gnd
rlabel metal1 2591 572 2595 573 1 Vdd
rlabel m2contact 2584 588 2588 592 7 Qbar
rlabel pdcontact 2571 588 2575 592 7 Dbar
rlabel m2contact 2584 577 2588 581 1 Q
rlabel pdcontact 2571 577 2575 581 1 D
rlabel polysilicon 2576 572 2578 573 1 En
rlabel polysilicon 2633 572 2635 573 1 En
rlabel metal1 2662 579 2666 583 7 Qout
rlabel pdcontact 2670 587 2674 591 7 Vdd
rlabel ndcontact 2654 587 2658 591 3 Gnd
rlabel metal1 2635 619 2639 620 6 Gnd
rlabel metal1 2591 596 2595 597 1 Vdd
rlabel m2contact 2584 612 2588 616 7 Qbar
rlabel pdcontact 2571 612 2575 616 7 Dbar
rlabel m2contact 2584 601 2588 605 1 Q
rlabel pdcontact 2571 601 2575 605 1 D
rlabel polysilicon 2576 596 2578 597 1 En
rlabel polysilicon 2633 596 2635 597 1 En
rlabel metal1 2662 603 2666 607 7 Qout
rlabel pdcontact 2670 611 2674 615 7 Vdd
rlabel ndcontact 2654 611 2658 615 3 Gnd
rlabel polysilicon 2484 644 2486 645 5 A
rlabel metal1 2483 636 2487 637 1 Z
rlabel metal1 2467 644 2471 645 4 Gnd
rlabel metal1 2499 644 2503 645 6 Vdd
rlabel metal1 2467 636 2471 637 8 Gnd
rlabel metal1 2435 636 2439 637 2 Vdd
rlabel polysilicon 2452 644 2454 645 5 A
rlabel metal1 2451 636 2455 637 1 Z
rlabel metal1 2515 595 2519 596 1 Gnd
rlabel metal1 2453 621 2456 622 5 Dbar
rlabel metal1 2388 595 2392 596 2 Gnd
rlabel metal1 2453 595 2456 596 1 Qbar
rlabel metal1 2460 595 2461 598 1 Q
rlabel polysilicon 2449 595 2451 596 1 Clk
rlabel metal1 2432 595 2436 596 1 Vdd
rlabel polysilicon 2557 621 2559 622 5 Clk
rlabel metal1 2559 595 2563 596 8 Vdd
rlabel polysilicon 2392 621 2394 622 5 Clk
rlabel metal1 2460 621 2463 622 5 D
rlabel polysilicon 2494 621 2502 622 5 En
rlabel polysilicon 2483 621 2491 622 5 Clk
rlabel metal1 2515 568 2519 569 1 Gnd
rlabel metal1 2453 594 2456 595 5 Dbar
rlabel metal1 2388 568 2392 569 2 Gnd
rlabel metal1 2453 568 2456 569 1 Qbar
rlabel metal1 2460 568 2461 571 1 Q
rlabel polysilicon 2449 568 2451 569 1 Clk
rlabel metal1 2432 568 2436 569 1 Vdd
rlabel polysilicon 2557 594 2559 595 5 Clk
rlabel metal1 2559 568 2563 569 8 Vdd
rlabel polysilicon 2392 594 2394 595 5 Clk
rlabel metal1 2460 594 2463 595 5 D
rlabel polysilicon 2494 594 2502 595 5 En
rlabel polysilicon 2483 594 2491 595 5 Clk
rlabel metal1 2515 541 2519 542 1 Gnd
rlabel metal1 2453 567 2456 568 5 Dbar
rlabel metal1 2388 541 2392 542 2 Gnd
rlabel metal1 2453 541 2456 542 1 Qbar
rlabel metal1 2460 541 2461 544 1 Q
rlabel polysilicon 2449 541 2451 542 1 Clk
rlabel metal1 2432 541 2436 542 1 Vdd
rlabel polysilicon 2557 567 2559 568 5 Clk
rlabel metal1 2559 541 2563 542 8 Vdd
rlabel polysilicon 2392 567 2394 568 5 Clk
rlabel metal1 2460 567 2463 568 5 D
rlabel polysilicon 2494 567 2502 568 5 En
rlabel polysilicon 2483 567 2491 568 5 Clk
rlabel metal1 2515 514 2519 515 1 Gnd
rlabel metal1 2453 540 2456 541 5 Dbar
rlabel metal1 2388 514 2392 515 2 Gnd
rlabel metal1 2453 514 2456 515 1 Qbar
rlabel metal1 2460 514 2461 517 1 Q
rlabel polysilicon 2449 514 2451 515 1 Clk
rlabel metal1 2432 514 2436 515 1 Vdd
rlabel polysilicon 2557 540 2559 541 5 Clk
rlabel metal1 2559 514 2563 515 8 Vdd
rlabel polysilicon 2392 540 2394 541 5 Clk
rlabel metal1 2460 540 2463 541 5 D
rlabel polysilicon 2494 540 2502 541 5 En
rlabel polysilicon 2483 540 2491 541 5 Clk
rlabel metal1 2860 4 2864 8 1 Gnd
rlabel metal1 2070 0 2074 4 1 Gnd
rlabel polysilicon 2758 526 2776 528 1 V+
rlabel polysilicon 2758 521 2776 523 1 V-
rlabel metal1 2690 520 2694 529 1 Gnd
rlabel metal1 2840 520 2844 529 1 Vdd
rlabel polysilicon 2738 398 2744 399 1 Vbp
rlabel polysilicon 2790 398 2796 399 1 Vbn
rlabel polysilicon 2821 398 2827 399 1 Vcp
rlabel polysilicon 2707 398 2713 399 1 Vcn
rlabel polysilicon 2695 398 2701 399 1 Vbn
rlabel polysilicon 2733 385 2739 387 5 Vbp
rlabel metal1 2692 253 2696 257 3 Vcn
rlabel metal1 2748 252 2752 264 1 Vbp
rlabel ndcontact 2740 241 2744 245 1 Gnd
rlabel pdcontact 2704 271 2708 275 1 Vdd
rlabel metal1 2784 252 2788 264 1 Vbn
rlabel metal1 2840 259 2844 263 7 Vcp
rlabel polysilicon 2797 129 2803 131 1 Vbn
rlabel ndcontact 2828 241 2832 245 1 Gnd
rlabel pdcontact 2792 271 2796 275 1 Vdd
rlabel ndcontact 2760 88 2764 92 1 M3source
rlabel ndcontact 2772 132 2776 136 1 Gnd
rlabel polysilicon 2753 384 2759 386 5 Vbp
rlabel pdiffusion 2783 382 2786 384 1 Vbn
rlabel pdiffusion 2839 382 2842 384 1 Vcp
rlabel polysilicon 2833 384 2839 386 5 Vcp
rlabel ndiffusion 2694 132 2697 134 1 Vcn
rlabel polysilicon 2697 130 2703 132 1 Vcn
rlabel pdiffusion 2694 382 2697 384 1 Vcn
<< end >>
