magic
tech scmos
timestamp 1418873681
<< end >>
