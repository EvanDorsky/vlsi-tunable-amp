magic
tech scmos
timestamp 1419285127
use bias  bias_0
timestamp 1418768461
transform 1 0 770 0 1 288
box 13 -282 183 102
use amp  amp_0
timestamp 1419283609
transform 1 0 781 0 1 394
box -781 -394 952 261
<< end >>
