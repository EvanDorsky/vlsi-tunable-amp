* SPICE3 file created from resistors.ext - technology: scmos

M1000 r1 c_5_n3# Vout Gnd phrResistor w=1.5u l=237.6u
+  ad=5.49p pd=10.2u as=4.14p ps=8.4u
M1001 r2 c_808_n3# r1 Gnd phrResistor w=1.5u l=15u
+  ad=5.04p pd=9.6u as=0p ps=0u
M1002 r3 c_868_n3# r2 Gnd phrResistor w=1.5u l=30u
+  ad=5.04p pd=9.6u as=0p ps=0u
M1003 r6 c_978_n3# r3 Gnd phrResistor w=1.5u l=15u
+  ad=5.04p pd=9.6u as=0p ps=0u
M1004 r4 c_1038_n3# r6 Gnd phrResistor w=1.5u l=60u
+  ad=5.04p pd=9.6u as=0p ps=0u
M1005 Vref c_1248_n3# r4 Gnd phrResistor w=1.5u l=120u
+  ad=4.14p pd=8.4u as=0p ps=0u
M1006 r2 B1 r3 Gnd nfet w=49.5u l=0.6u
+  ad=93.06p pd=208.2u as=45.27p ps=102u
M1007 r2 B0 r1 Gnd nfet w=49.5u l=0.6u
+  ad=0p pd=0u as=45.27p ps=102u
M1008 r6 B2 r4 Gnd nfet w=49.5u l=0.6u
+  ad=45.27p pd=102u as=90.54p ps=204u
M1009 r4 B3 Vref Gnd nfet w=49.5u l=0.6u
+  ad=0p pd=0u as=45.27p ps=102u
C0 r1 r3 3.8fF
