magic
tech scmos
timestamp 1417655414
<< ntransistor >>
rect -5 -18 -1 -16
rect 6 -18 10 -16
rect -7 -44 -4 -38
rect 0 -44 3 -38
rect -5 -123 -1 -121
rect 6 -123 10 -121
rect 0 -130 5 -128
<< ptransistor >>
rect 0 19 5 21
rect -5 12 -1 14
rect 6 12 10 14
rect -8 -71 -4 -69
rect 0 -71 4 -69
rect -5 -93 -1 -91
rect 6 -93 10 -91
<< ndiffusion >>
rect -5 -16 -1 -15
rect 6 -16 10 -15
rect -5 -21 -1 -18
rect 6 -21 10 -18
rect -7 -38 -4 -37
rect 0 -38 3 -37
rect -7 -45 -4 -44
rect 0 -45 3 -44
rect -5 -121 -1 -120
rect 6 -121 10 -120
rect -5 -124 -1 -123
rect 6 -124 10 -123
rect -5 -127 10 -124
rect 0 -128 5 -127
rect 0 -131 5 -130
rect -1 -134 6 -131
<< pdiffusion >>
rect -1 22 6 25
rect 0 21 5 22
rect 0 18 5 19
rect -5 15 10 18
rect -5 14 -1 15
rect 6 14 10 15
rect -5 11 -1 12
rect 6 11 10 12
rect -8 -69 -4 -68
rect 0 -69 4 -68
rect -8 -72 -4 -71
rect 0 -72 4 -71
rect -5 -91 -1 -88
rect 6 -91 10 -88
rect -5 -94 -1 -93
rect 6 -94 10 -93
<< ndcontact >>
rect -5 -15 -1 -11
rect 6 -15 10 -11
rect -5 -25 -1 -21
rect 6 -25 10 -21
rect -8 -37 -4 -33
rect 0 -37 4 -33
rect -8 -49 -4 -45
rect 0 -49 4 -45
rect -5 -120 -1 -116
rect 6 -120 10 -116
rect -5 -135 -1 -131
rect 6 -135 10 -131
<< pdcontact >>
rect -5 22 -1 26
rect 6 22 10 26
rect -5 7 -1 11
rect 6 7 10 11
rect -8 -68 -4 -64
rect 0 -68 4 -64
rect -8 -76 -4 -72
rect 0 -76 4 -72
rect -5 -88 -1 -84
rect 6 -88 10 -84
rect -5 -98 -1 -94
rect 6 -98 10 -94
<< polysilicon >>
rect -11 19 0 21
rect 5 19 16 21
rect -8 12 -5 14
rect -1 12 1 14
rect 4 12 6 14
rect 10 12 13 14
rect -8 -6 -6 12
rect 11 4 13 12
rect 3 2 13 4
rect -8 -8 2 -6
rect -8 -16 -6 -8
rect 11 -16 13 2
rect -8 -18 -5 -16
rect -1 -18 1 -16
rect 4 -18 6 -16
rect 10 -18 13 -16
rect -11 -44 -7 -38
rect -4 -44 0 -38
rect 3 -44 16 -38
rect -11 -71 -8 -69
rect -4 -71 0 -69
rect 4 -71 16 -69
rect -8 -93 -5 -91
rect -1 -93 1 -91
rect 4 -93 6 -91
rect 10 -93 13 -91
rect -8 -111 -6 -93
rect 11 -101 13 -93
rect 3 -103 13 -101
rect -8 -113 2 -111
rect -8 -121 -6 -113
rect 11 -121 13 -103
rect -8 -123 -5 -121
rect -1 -123 1 -121
rect 4 -123 6 -121
rect 10 -123 13 -121
rect -11 -130 0 -128
rect 5 -130 16 -128
<< polycontact >>
rect -1 1 3 5
rect 2 -9 6 -5
rect -1 -104 3 -100
rect 2 -114 6 -110
<< metal1 >>
rect -11 22 -5 25
rect -1 22 6 25
rect 10 22 16 25
rect -11 21 16 22
rect -5 0 -1 7
rect -5 -11 -1 -4
rect 6 0 10 7
rect 6 -11 10 -4
rect -11 -25 -5 -21
rect -1 -25 6 -21
rect 10 -25 16 -21
rect -8 -33 -4 -32
rect 0 -33 4 -32
rect -8 -50 -4 -49
rect 0 -50 3 -49
rect 7 -51 10 -38
rect 7 -54 16 -51
rect -11 -60 2 -57
rect -1 -64 2 -60
rect 13 -60 16 -54
rect 7 -64 10 -61
rect -1 -68 0 -64
rect 7 -67 16 -64
rect -8 -77 -4 -76
rect 0 -77 4 -76
rect -11 -88 -5 -84
rect -1 -88 6 -84
rect 10 -88 16 -84
rect -5 -105 -1 -98
rect -5 -116 -1 -109
rect 6 -105 10 -98
rect 6 -116 10 -109
rect -11 -131 16 -130
rect -11 -134 -5 -131
rect -1 -134 6 -131
rect 10 -134 16 -131
<< m2contact >>
rect -5 -4 -1 0
rect 6 -4 10 0
rect -8 -32 -4 -28
rect 0 -32 4 -28
rect 7 -38 11 -34
rect -8 -54 -4 -50
rect -1 -54 3 -50
rect 6 -61 10 -57
rect -8 -81 -4 -77
rect 0 -81 4 -77
rect -5 -109 -1 -105
rect 6 -109 10 -105
<< metal2 >>
rect -5 -18 -1 -4
rect -8 -21 -1 -18
rect -8 -28 -4 -21
rect 6 -25 10 -4
rect 0 -28 10 -25
rect -7 -42 -4 -32
rect 7 -34 10 -28
rect -7 -45 9 -42
rect -8 -77 -5 -54
rect -1 -77 2 -54
rect 6 -57 9 -45
rect -1 -81 0 -77
rect -8 -109 -5 -81
rect -1 -105 2 -81
rect -1 -109 6 -105
<< labels >>
rlabel pdcontact -5 -68 -4 -64 1 Dbar
rlabel metal1 -5 -60 -4 -57 1 D
rlabel polysilicon -8 -44 -7 -38 3 Clk
rlabel polysilicon -8 19 -7 21 3 Clk
rlabel metal1 -8 21 -7 25 4 Vdd
rlabel metal1 15 -88 16 -84 7 Vdd
rlabel polysilicon 15 -71 16 -69 7 Clk
rlabel metal1 13 -60 16 -59 7 Q
rlabel metal1 15 -67 16 -64 7 Qbar
rlabel metal1 15 -25 16 -21 7 Gnd
rlabel metal1 15 -134 16 -130 8 Gnd
rlabel polysilicon -8 -130 -7 -128 3 Clk
<< end >>
