magic
tech scmos
timestamp 1259953556
<< electrodecontact >>
rect 384 4090 388 4094
rect 397 4090 401 4094
rect 384 4084 388 4088
rect 397 4084 401 4088
rect 384 4078 388 4082
rect 397 4078 401 4082
rect 384 4072 388 4076
rect 397 4072 401 4076
rect 384 4066 388 4070
rect 397 4066 401 4070
rect 414 4089 418 4093
rect 420 4089 424 4093
rect 427 4089 431 4093
rect 433 4089 437 4093
rect 439 4089 443 4093
rect 445 4089 449 4093
rect 471 4090 475 4094
rect 489 4090 493 4094
rect 414 4083 418 4087
rect 420 4083 424 4087
rect 427 4083 431 4087
rect 433 4083 437 4087
rect 439 4083 443 4087
rect 445 4083 449 4087
rect 471 4084 475 4088
rect 489 4084 493 4088
rect 414 4077 418 4081
rect 420 4077 424 4081
rect 427 4077 431 4081
rect 433 4077 437 4081
rect 439 4077 443 4081
rect 445 4077 449 4081
rect 471 4078 475 4082
rect 489 4078 493 4082
rect 414 4071 418 4075
rect 420 4071 424 4075
rect 427 4071 431 4075
rect 433 4071 437 4075
rect 439 4071 443 4075
rect 445 4071 449 4075
rect 471 4072 475 4076
rect 489 4072 493 4076
rect 414 4065 418 4069
rect 420 4065 424 4069
rect 427 4065 431 4069
rect 433 4065 437 4069
rect 439 4065 443 4069
rect 445 4065 449 4069
rect 471 4066 475 4070
rect 489 4066 493 4070
rect 384 4060 388 4064
rect 397 4060 401 4064
rect 471 4060 475 4064
rect 489 4060 493 4064
rect 384 4054 388 4058
rect 397 4054 401 4058
rect 456 4056 460 4060
rect 471 4054 475 4058
rect 489 4054 493 4058
rect 456 4046 460 4050
rect 456 4008 460 4012
rect 384 4000 388 4004
rect 397 4000 401 4004
rect 456 3998 460 4002
rect 471 4000 475 4004
rect 489 4000 493 4004
rect 384 3994 388 3998
rect 397 3994 401 3998
rect 471 3994 475 3998
rect 489 3994 493 3998
rect 384 3988 388 3992
rect 397 3988 401 3992
rect 384 3982 388 3986
rect 397 3982 401 3986
rect 384 3976 388 3980
rect 397 3976 401 3980
rect 384 3970 388 3974
rect 397 3970 401 3974
rect 384 3964 388 3968
rect 397 3964 401 3968
rect 414 3989 418 3993
rect 420 3989 424 3993
rect 427 3989 431 3993
rect 433 3989 437 3993
rect 439 3989 443 3993
rect 445 3989 449 3993
rect 471 3988 475 3992
rect 489 3988 493 3992
rect 414 3983 418 3987
rect 420 3983 424 3987
rect 427 3983 431 3987
rect 433 3983 437 3987
rect 439 3983 443 3987
rect 445 3983 449 3987
rect 471 3982 475 3986
rect 489 3982 493 3986
rect 414 3977 418 3981
rect 420 3977 424 3981
rect 427 3977 431 3981
rect 433 3977 437 3981
rect 439 3977 443 3981
rect 445 3977 449 3981
rect 471 3976 475 3980
rect 489 3976 493 3980
rect 414 3971 418 3975
rect 420 3971 424 3975
rect 427 3971 431 3975
rect 433 3971 437 3975
rect 439 3971 443 3975
rect 445 3971 449 3975
rect 471 3970 475 3974
rect 489 3970 493 3974
rect 414 3965 418 3969
rect 420 3965 424 3969
rect 427 3965 431 3969
rect 433 3965 437 3969
rect 439 3965 443 3969
rect 445 3965 449 3969
rect 471 3964 475 3968
rect 489 3964 493 3968
rect 384 3616 388 3620
rect 397 3616 401 3620
rect 384 3610 388 3614
rect 397 3610 401 3614
rect 384 3604 388 3608
rect 397 3604 401 3608
rect 384 3598 388 3602
rect 397 3598 401 3602
rect 384 3592 388 3596
rect 397 3592 401 3596
rect 414 3615 418 3619
rect 420 3615 424 3619
rect 427 3615 431 3619
rect 433 3615 437 3619
rect 439 3615 443 3619
rect 445 3615 449 3619
rect 471 3616 475 3620
rect 489 3616 493 3620
rect 414 3609 418 3613
rect 420 3609 424 3613
rect 427 3609 431 3613
rect 433 3609 437 3613
rect 439 3609 443 3613
rect 445 3609 449 3613
rect 471 3610 475 3614
rect 489 3610 493 3614
rect 414 3603 418 3607
rect 420 3603 424 3607
rect 427 3603 431 3607
rect 433 3603 437 3607
rect 439 3603 443 3607
rect 445 3603 449 3607
rect 471 3604 475 3608
rect 489 3604 493 3608
rect 414 3597 418 3601
rect 420 3597 424 3601
rect 427 3597 431 3601
rect 433 3597 437 3601
rect 439 3597 443 3601
rect 445 3597 449 3601
rect 471 3598 475 3602
rect 489 3598 493 3602
rect 414 3591 418 3595
rect 420 3591 424 3595
rect 427 3591 431 3595
rect 433 3591 437 3595
rect 439 3591 443 3595
rect 445 3591 449 3595
rect 471 3592 475 3596
rect 489 3592 493 3596
rect 384 3586 388 3590
rect 397 3586 401 3590
rect 471 3586 475 3590
rect 489 3586 493 3590
rect 384 3580 388 3584
rect 397 3580 401 3584
rect 456 3582 460 3586
rect 471 3580 475 3584
rect 489 3580 493 3584
rect 456 3572 460 3576
rect 456 3534 460 3538
rect 384 3526 388 3530
rect 397 3526 401 3530
rect 456 3524 460 3528
rect 471 3526 475 3530
rect 489 3526 493 3530
rect 384 3520 388 3524
rect 397 3520 401 3524
rect 471 3520 475 3524
rect 489 3520 493 3524
rect 384 3514 388 3518
rect 397 3514 401 3518
rect 384 3508 388 3512
rect 397 3508 401 3512
rect 384 3502 388 3506
rect 397 3502 401 3506
rect 384 3496 388 3500
rect 397 3496 401 3500
rect 384 3490 388 3494
rect 397 3490 401 3494
rect 414 3515 418 3519
rect 420 3515 424 3519
rect 427 3515 431 3519
rect 433 3515 437 3519
rect 439 3515 443 3519
rect 445 3515 449 3519
rect 471 3514 475 3518
rect 489 3514 493 3518
rect 414 3509 418 3513
rect 420 3509 424 3513
rect 427 3509 431 3513
rect 433 3509 437 3513
rect 439 3509 443 3513
rect 445 3509 449 3513
rect 471 3508 475 3512
rect 489 3508 493 3512
rect 414 3503 418 3507
rect 420 3503 424 3507
rect 427 3503 431 3507
rect 433 3503 437 3507
rect 439 3503 443 3507
rect 445 3503 449 3507
rect 471 3502 475 3506
rect 489 3502 493 3506
rect 414 3497 418 3501
rect 420 3497 424 3501
rect 427 3497 431 3501
rect 433 3497 437 3501
rect 439 3497 443 3501
rect 445 3497 449 3501
rect 471 3496 475 3500
rect 489 3496 493 3500
rect 414 3491 418 3495
rect 420 3491 424 3495
rect 427 3491 431 3495
rect 433 3491 437 3495
rect 439 3491 443 3495
rect 445 3491 449 3495
rect 471 3490 475 3494
rect 489 3490 493 3494
rect 384 3142 388 3146
rect 397 3142 401 3146
rect 384 3136 388 3140
rect 397 3136 401 3140
rect 384 3130 388 3134
rect 397 3130 401 3134
rect 384 3124 388 3128
rect 397 3124 401 3128
rect 384 3118 388 3122
rect 397 3118 401 3122
rect 414 3141 418 3145
rect 420 3141 424 3145
rect 427 3141 431 3145
rect 433 3141 437 3145
rect 439 3141 443 3145
rect 445 3141 449 3145
rect 471 3142 475 3146
rect 489 3142 493 3146
rect 414 3135 418 3139
rect 420 3135 424 3139
rect 427 3135 431 3139
rect 433 3135 437 3139
rect 439 3135 443 3139
rect 445 3135 449 3139
rect 471 3136 475 3140
rect 489 3136 493 3140
rect 414 3129 418 3133
rect 420 3129 424 3133
rect 427 3129 431 3133
rect 433 3129 437 3133
rect 439 3129 443 3133
rect 445 3129 449 3133
rect 471 3130 475 3134
rect 489 3130 493 3134
rect 414 3123 418 3127
rect 420 3123 424 3127
rect 427 3123 431 3127
rect 433 3123 437 3127
rect 439 3123 443 3127
rect 445 3123 449 3127
rect 471 3124 475 3128
rect 489 3124 493 3128
rect 414 3117 418 3121
rect 420 3117 424 3121
rect 427 3117 431 3121
rect 433 3117 437 3121
rect 439 3117 443 3121
rect 445 3117 449 3121
rect 471 3118 475 3122
rect 489 3118 493 3122
rect 384 3112 388 3116
rect 397 3112 401 3116
rect 471 3112 475 3116
rect 489 3112 493 3116
rect 384 3106 388 3110
rect 397 3106 401 3110
rect 456 3108 460 3112
rect 471 3106 475 3110
rect 489 3106 493 3110
rect 456 3098 460 3102
rect 456 3060 460 3064
rect 384 3052 388 3056
rect 397 3052 401 3056
rect 456 3050 460 3054
rect 471 3052 475 3056
rect 489 3052 493 3056
rect 384 3046 388 3050
rect 397 3046 401 3050
rect 471 3046 475 3050
rect 489 3046 493 3050
rect 384 3040 388 3044
rect 397 3040 401 3044
rect 384 3034 388 3038
rect 397 3034 401 3038
rect 384 3028 388 3032
rect 397 3028 401 3032
rect 384 3022 388 3026
rect 397 3022 401 3026
rect 384 3016 388 3020
rect 397 3016 401 3020
rect 414 3041 418 3045
rect 420 3041 424 3045
rect 427 3041 431 3045
rect 433 3041 437 3045
rect 439 3041 443 3045
rect 445 3041 449 3045
rect 471 3040 475 3044
rect 489 3040 493 3044
rect 414 3035 418 3039
rect 420 3035 424 3039
rect 427 3035 431 3039
rect 433 3035 437 3039
rect 439 3035 443 3039
rect 445 3035 449 3039
rect 471 3034 475 3038
rect 489 3034 493 3038
rect 414 3029 418 3033
rect 420 3029 424 3033
rect 427 3029 431 3033
rect 433 3029 437 3033
rect 439 3029 443 3033
rect 445 3029 449 3033
rect 471 3028 475 3032
rect 489 3028 493 3032
rect 414 3023 418 3027
rect 420 3023 424 3027
rect 427 3023 431 3027
rect 433 3023 437 3027
rect 439 3023 443 3027
rect 445 3023 449 3027
rect 471 3022 475 3026
rect 489 3022 493 3026
rect 414 3017 418 3021
rect 420 3017 424 3021
rect 427 3017 431 3021
rect 433 3017 437 3021
rect 439 3017 443 3021
rect 445 3017 449 3021
rect 471 3016 475 3020
rect 489 3016 493 3020
rect 384 2668 388 2672
rect 397 2668 401 2672
rect 384 2662 388 2666
rect 397 2662 401 2666
rect 384 2656 388 2660
rect 397 2656 401 2660
rect 384 2650 388 2654
rect 397 2650 401 2654
rect 384 2644 388 2648
rect 397 2644 401 2648
rect 414 2667 418 2671
rect 420 2667 424 2671
rect 427 2667 431 2671
rect 433 2667 437 2671
rect 439 2667 443 2671
rect 445 2667 449 2671
rect 471 2668 475 2672
rect 489 2668 493 2672
rect 414 2661 418 2665
rect 420 2661 424 2665
rect 427 2661 431 2665
rect 433 2661 437 2665
rect 439 2661 443 2665
rect 445 2661 449 2665
rect 471 2662 475 2666
rect 489 2662 493 2666
rect 414 2655 418 2659
rect 420 2655 424 2659
rect 427 2655 431 2659
rect 433 2655 437 2659
rect 439 2655 443 2659
rect 445 2655 449 2659
rect 471 2656 475 2660
rect 489 2656 493 2660
rect 414 2649 418 2653
rect 420 2649 424 2653
rect 427 2649 431 2653
rect 433 2649 437 2653
rect 439 2649 443 2653
rect 445 2649 449 2653
rect 471 2650 475 2654
rect 489 2650 493 2654
rect 414 2643 418 2647
rect 420 2643 424 2647
rect 427 2643 431 2647
rect 433 2643 437 2647
rect 439 2643 443 2647
rect 445 2643 449 2647
rect 471 2644 475 2648
rect 489 2644 493 2648
rect 384 2638 388 2642
rect 397 2638 401 2642
rect 471 2638 475 2642
rect 489 2638 493 2642
rect 384 2632 388 2636
rect 397 2632 401 2636
rect 456 2634 460 2638
rect 471 2632 475 2636
rect 489 2632 493 2636
rect 456 2624 460 2628
rect 456 2586 460 2590
rect 384 2578 388 2582
rect 397 2578 401 2582
rect 456 2576 460 2580
rect 471 2578 475 2582
rect 489 2578 493 2582
rect 384 2572 388 2576
rect 397 2572 401 2576
rect 471 2572 475 2576
rect 489 2572 493 2576
rect 384 2566 388 2570
rect 397 2566 401 2570
rect 384 2560 388 2564
rect 397 2560 401 2564
rect 384 2554 388 2558
rect 397 2554 401 2558
rect 384 2548 388 2552
rect 397 2548 401 2552
rect 384 2542 388 2546
rect 397 2542 401 2546
rect 414 2567 418 2571
rect 420 2567 424 2571
rect 427 2567 431 2571
rect 433 2567 437 2571
rect 439 2567 443 2571
rect 445 2567 449 2571
rect 471 2566 475 2570
rect 489 2566 493 2570
rect 414 2561 418 2565
rect 420 2561 424 2565
rect 427 2561 431 2565
rect 433 2561 437 2565
rect 439 2561 443 2565
rect 445 2561 449 2565
rect 471 2560 475 2564
rect 489 2560 493 2564
rect 414 2555 418 2559
rect 420 2555 424 2559
rect 427 2555 431 2559
rect 433 2555 437 2559
rect 439 2555 443 2559
rect 445 2555 449 2559
rect 471 2554 475 2558
rect 489 2554 493 2558
rect 414 2549 418 2553
rect 420 2549 424 2553
rect 427 2549 431 2553
rect 433 2549 437 2553
rect 439 2549 443 2553
rect 445 2549 449 2553
rect 471 2548 475 2552
rect 489 2548 493 2552
rect 414 2543 418 2547
rect 420 2543 424 2547
rect 427 2543 431 2547
rect 433 2543 437 2547
rect 439 2543 443 2547
rect 445 2543 449 2547
rect 471 2542 475 2546
rect 489 2542 493 2546
rect 384 2194 388 2198
rect 397 2194 401 2198
rect 384 2188 388 2192
rect 397 2188 401 2192
rect 384 2182 388 2186
rect 397 2182 401 2186
rect 384 2176 388 2180
rect 397 2176 401 2180
rect 384 2170 388 2174
rect 397 2170 401 2174
rect 414 2193 418 2197
rect 420 2193 424 2197
rect 427 2193 431 2197
rect 433 2193 437 2197
rect 439 2193 443 2197
rect 445 2193 449 2197
rect 471 2194 475 2198
rect 489 2194 493 2198
rect 414 2187 418 2191
rect 420 2187 424 2191
rect 427 2187 431 2191
rect 433 2187 437 2191
rect 439 2187 443 2191
rect 445 2187 449 2191
rect 471 2188 475 2192
rect 489 2188 493 2192
rect 414 2181 418 2185
rect 420 2181 424 2185
rect 427 2181 431 2185
rect 433 2181 437 2185
rect 439 2181 443 2185
rect 445 2181 449 2185
rect 471 2182 475 2186
rect 489 2182 493 2186
rect 414 2175 418 2179
rect 420 2175 424 2179
rect 427 2175 431 2179
rect 433 2175 437 2179
rect 439 2175 443 2179
rect 445 2175 449 2179
rect 471 2176 475 2180
rect 489 2176 493 2180
rect 414 2169 418 2173
rect 420 2169 424 2173
rect 427 2169 431 2173
rect 433 2169 437 2173
rect 439 2169 443 2173
rect 445 2169 449 2173
rect 471 2170 475 2174
rect 489 2170 493 2174
rect 384 2164 388 2168
rect 397 2164 401 2168
rect 471 2164 475 2168
rect 489 2164 493 2168
rect 384 2158 388 2162
rect 397 2158 401 2162
rect 456 2160 460 2164
rect 471 2158 475 2162
rect 489 2158 493 2162
rect 456 2150 460 2154
rect 456 2112 460 2116
rect 384 2104 388 2108
rect 397 2104 401 2108
rect 456 2102 460 2106
rect 471 2104 475 2108
rect 489 2104 493 2108
rect 384 2098 388 2102
rect 397 2098 401 2102
rect 471 2098 475 2102
rect 489 2098 493 2102
rect 384 2092 388 2096
rect 397 2092 401 2096
rect 384 2086 388 2090
rect 397 2086 401 2090
rect 384 2080 388 2084
rect 397 2080 401 2084
rect 384 2074 388 2078
rect 397 2074 401 2078
rect 384 2068 388 2072
rect 397 2068 401 2072
rect 414 2093 418 2097
rect 420 2093 424 2097
rect 427 2093 431 2097
rect 433 2093 437 2097
rect 439 2093 443 2097
rect 445 2093 449 2097
rect 471 2092 475 2096
rect 489 2092 493 2096
rect 414 2087 418 2091
rect 420 2087 424 2091
rect 427 2087 431 2091
rect 433 2087 437 2091
rect 439 2087 443 2091
rect 445 2087 449 2091
rect 471 2086 475 2090
rect 489 2086 493 2090
rect 414 2081 418 2085
rect 420 2081 424 2085
rect 427 2081 431 2085
rect 433 2081 437 2085
rect 439 2081 443 2085
rect 445 2081 449 2085
rect 471 2080 475 2084
rect 489 2080 493 2084
rect 414 2075 418 2079
rect 420 2075 424 2079
rect 427 2075 431 2079
rect 433 2075 437 2079
rect 439 2075 443 2079
rect 445 2075 449 2079
rect 471 2074 475 2078
rect 489 2074 493 2078
rect 414 2069 418 2073
rect 420 2069 424 2073
rect 427 2069 431 2073
rect 433 2069 437 2073
rect 439 2069 443 2073
rect 445 2069 449 2073
rect 471 2068 475 2072
rect 489 2068 493 2072
rect 384 1720 388 1724
rect 397 1720 401 1724
rect 384 1714 388 1718
rect 397 1714 401 1718
rect 384 1708 388 1712
rect 397 1708 401 1712
rect 384 1702 388 1706
rect 397 1702 401 1706
rect 384 1696 388 1700
rect 397 1696 401 1700
rect 414 1719 418 1723
rect 420 1719 424 1723
rect 427 1719 431 1723
rect 433 1719 437 1723
rect 439 1719 443 1723
rect 445 1719 449 1723
rect 471 1720 475 1724
rect 489 1720 493 1724
rect 414 1713 418 1717
rect 420 1713 424 1717
rect 427 1713 431 1717
rect 433 1713 437 1717
rect 439 1713 443 1717
rect 445 1713 449 1717
rect 471 1714 475 1718
rect 489 1714 493 1718
rect 414 1707 418 1711
rect 420 1707 424 1711
rect 427 1707 431 1711
rect 433 1707 437 1711
rect 439 1707 443 1711
rect 445 1707 449 1711
rect 471 1708 475 1712
rect 489 1708 493 1712
rect 414 1701 418 1705
rect 420 1701 424 1705
rect 427 1701 431 1705
rect 433 1701 437 1705
rect 439 1701 443 1705
rect 445 1701 449 1705
rect 471 1702 475 1706
rect 489 1702 493 1706
rect 414 1695 418 1699
rect 420 1695 424 1699
rect 427 1695 431 1699
rect 433 1695 437 1699
rect 439 1695 443 1699
rect 445 1695 449 1699
rect 471 1696 475 1700
rect 489 1696 493 1700
rect 384 1690 388 1694
rect 397 1690 401 1694
rect 471 1690 475 1694
rect 489 1690 493 1694
rect 384 1684 388 1688
rect 397 1684 401 1688
rect 456 1686 460 1690
rect 471 1684 475 1688
rect 489 1684 493 1688
rect 456 1676 460 1680
rect 456 1638 460 1642
rect 384 1630 388 1634
rect 397 1630 401 1634
rect 456 1628 460 1632
rect 471 1630 475 1634
rect 489 1630 493 1634
rect 384 1624 388 1628
rect 397 1624 401 1628
rect 471 1624 475 1628
rect 489 1624 493 1628
rect 384 1618 388 1622
rect 397 1618 401 1622
rect 384 1612 388 1616
rect 397 1612 401 1616
rect 384 1606 388 1610
rect 397 1606 401 1610
rect 384 1600 388 1604
rect 397 1600 401 1604
rect 384 1594 388 1598
rect 397 1594 401 1598
rect 414 1619 418 1623
rect 420 1619 424 1623
rect 427 1619 431 1623
rect 433 1619 437 1623
rect 439 1619 443 1623
rect 445 1619 449 1623
rect 471 1618 475 1622
rect 489 1618 493 1622
rect 414 1613 418 1617
rect 420 1613 424 1617
rect 427 1613 431 1617
rect 433 1613 437 1617
rect 439 1613 443 1617
rect 445 1613 449 1617
rect 471 1612 475 1616
rect 489 1612 493 1616
rect 414 1607 418 1611
rect 420 1607 424 1611
rect 427 1607 431 1611
rect 433 1607 437 1611
rect 439 1607 443 1611
rect 445 1607 449 1611
rect 471 1606 475 1610
rect 489 1606 493 1610
rect 414 1601 418 1605
rect 420 1601 424 1605
rect 427 1601 431 1605
rect 433 1601 437 1605
rect 439 1601 443 1605
rect 445 1601 449 1605
rect 471 1600 475 1604
rect 489 1600 493 1604
rect 414 1595 418 1599
rect 420 1595 424 1599
rect 427 1595 431 1599
rect 433 1595 437 1599
rect 439 1595 443 1599
rect 445 1595 449 1599
rect 471 1594 475 1598
rect 489 1594 493 1598
rect 384 1246 388 1250
rect 397 1246 401 1250
rect 384 1240 388 1244
rect 397 1240 401 1244
rect 384 1234 388 1238
rect 397 1234 401 1238
rect 384 1228 388 1232
rect 397 1228 401 1232
rect 384 1222 388 1226
rect 397 1222 401 1226
rect 414 1245 418 1249
rect 420 1245 424 1249
rect 427 1245 431 1249
rect 433 1245 437 1249
rect 439 1245 443 1249
rect 445 1245 449 1249
rect 471 1246 475 1250
rect 489 1246 493 1250
rect 414 1239 418 1243
rect 420 1239 424 1243
rect 427 1239 431 1243
rect 433 1239 437 1243
rect 439 1239 443 1243
rect 445 1239 449 1243
rect 471 1240 475 1244
rect 489 1240 493 1244
rect 414 1233 418 1237
rect 420 1233 424 1237
rect 427 1233 431 1237
rect 433 1233 437 1237
rect 439 1233 443 1237
rect 445 1233 449 1237
rect 471 1234 475 1238
rect 489 1234 493 1238
rect 414 1227 418 1231
rect 420 1227 424 1231
rect 427 1227 431 1231
rect 433 1227 437 1231
rect 439 1227 443 1231
rect 445 1227 449 1231
rect 471 1228 475 1232
rect 489 1228 493 1232
rect 414 1221 418 1225
rect 420 1221 424 1225
rect 427 1221 431 1225
rect 433 1221 437 1225
rect 439 1221 443 1225
rect 445 1221 449 1225
rect 471 1222 475 1226
rect 489 1222 493 1226
rect 384 1216 388 1220
rect 397 1216 401 1220
rect 471 1216 475 1220
rect 489 1216 493 1220
rect 384 1210 388 1214
rect 397 1210 401 1214
rect 456 1212 460 1216
rect 471 1210 475 1214
rect 489 1210 493 1214
rect 456 1202 460 1206
rect 456 1164 460 1168
rect 384 1156 388 1160
rect 397 1156 401 1160
rect 456 1154 460 1158
rect 471 1156 475 1160
rect 489 1156 493 1160
rect 384 1150 388 1154
rect 397 1150 401 1154
rect 471 1150 475 1154
rect 489 1150 493 1154
rect 384 1144 388 1148
rect 397 1144 401 1148
rect 384 1138 388 1142
rect 397 1138 401 1142
rect 384 1132 388 1136
rect 397 1132 401 1136
rect 384 1126 388 1130
rect 397 1126 401 1130
rect 384 1120 388 1124
rect 397 1120 401 1124
rect 414 1145 418 1149
rect 420 1145 424 1149
rect 427 1145 431 1149
rect 433 1145 437 1149
rect 439 1145 443 1149
rect 445 1145 449 1149
rect 471 1144 475 1148
rect 489 1144 493 1148
rect 414 1139 418 1143
rect 420 1139 424 1143
rect 427 1139 431 1143
rect 433 1139 437 1143
rect 439 1139 443 1143
rect 445 1139 449 1143
rect 471 1138 475 1142
rect 489 1138 493 1142
rect 414 1133 418 1137
rect 420 1133 424 1137
rect 427 1133 431 1137
rect 433 1133 437 1137
rect 439 1133 443 1137
rect 445 1133 449 1137
rect 471 1132 475 1136
rect 489 1132 493 1136
rect 414 1127 418 1131
rect 420 1127 424 1131
rect 427 1127 431 1131
rect 433 1127 437 1131
rect 439 1127 443 1131
rect 445 1127 449 1131
rect 471 1126 475 1130
rect 489 1126 493 1130
rect 414 1121 418 1125
rect 420 1121 424 1125
rect 427 1121 431 1125
rect 433 1121 437 1125
rect 439 1121 443 1125
rect 445 1121 449 1125
rect 471 1120 475 1124
rect 489 1120 493 1124
rect 384 772 388 776
rect 397 772 401 776
rect 384 766 388 770
rect 397 766 401 770
rect 384 760 388 764
rect 397 760 401 764
rect 384 754 388 758
rect 397 754 401 758
rect 384 748 388 752
rect 397 748 401 752
rect 414 771 418 775
rect 420 771 424 775
rect 427 771 431 775
rect 433 771 437 775
rect 439 771 443 775
rect 445 771 449 775
rect 471 772 475 776
rect 489 772 493 776
rect 414 765 418 769
rect 420 765 424 769
rect 427 765 431 769
rect 433 765 437 769
rect 439 765 443 769
rect 445 765 449 769
rect 471 766 475 770
rect 489 766 493 770
rect 414 759 418 763
rect 420 759 424 763
rect 427 759 431 763
rect 433 759 437 763
rect 439 759 443 763
rect 445 759 449 763
rect 471 760 475 764
rect 489 760 493 764
rect 414 753 418 757
rect 420 753 424 757
rect 427 753 431 757
rect 433 753 437 757
rect 439 753 443 757
rect 445 753 449 757
rect 471 754 475 758
rect 489 754 493 758
rect 414 747 418 751
rect 420 747 424 751
rect 427 747 431 751
rect 433 747 437 751
rect 439 747 443 751
rect 445 747 449 751
rect 471 748 475 752
rect 489 748 493 752
rect 384 742 388 746
rect 397 742 401 746
rect 471 742 475 746
rect 489 742 493 746
rect 384 736 388 740
rect 397 736 401 740
rect 456 738 460 742
rect 471 736 475 740
rect 489 736 493 740
rect 456 728 460 732
rect 456 690 460 694
rect 384 682 388 686
rect 397 682 401 686
rect 456 680 460 684
rect 471 682 475 686
rect 489 682 493 686
rect 384 676 388 680
rect 397 676 401 680
rect 471 676 475 680
rect 489 676 493 680
rect 384 670 388 674
rect 397 670 401 674
rect 384 664 388 668
rect 397 664 401 668
rect 384 658 388 662
rect 397 658 401 662
rect 384 652 388 656
rect 397 652 401 656
rect 384 646 388 650
rect 397 646 401 650
rect 414 671 418 675
rect 420 671 424 675
rect 427 671 431 675
rect 433 671 437 675
rect 439 671 443 675
rect 445 671 449 675
rect 471 670 475 674
rect 489 670 493 674
rect 414 665 418 669
rect 420 665 424 669
rect 427 665 431 669
rect 433 665 437 669
rect 439 665 443 669
rect 445 665 449 669
rect 471 664 475 668
rect 489 664 493 668
rect 414 659 418 663
rect 420 659 424 663
rect 427 659 431 663
rect 433 659 437 663
rect 439 659 443 663
rect 445 659 449 663
rect 471 658 475 662
rect 489 658 493 662
rect 414 653 418 657
rect 420 653 424 657
rect 427 653 431 657
rect 433 653 437 657
rect 439 653 443 657
rect 445 653 449 657
rect 471 652 475 656
rect 489 652 493 656
rect 414 647 418 651
rect 420 647 424 651
rect 427 647 431 651
rect 433 647 437 651
rect 439 647 443 651
rect 445 647 449 651
rect 471 646 475 650
rect 489 646 493 650
rect 384 298 388 302
rect 397 298 401 302
rect 384 292 388 296
rect 397 292 401 296
rect 384 286 388 290
rect 397 286 401 290
rect 384 280 388 284
rect 397 280 401 284
rect 384 274 388 278
rect 397 274 401 278
rect 414 297 418 301
rect 420 297 424 301
rect 427 297 431 301
rect 433 297 437 301
rect 439 297 443 301
rect 445 297 449 301
rect 471 298 475 302
rect 489 298 493 302
rect 414 291 418 295
rect 420 291 424 295
rect 427 291 431 295
rect 433 291 437 295
rect 439 291 443 295
rect 445 291 449 295
rect 471 292 475 296
rect 489 292 493 296
rect 414 285 418 289
rect 420 285 424 289
rect 427 285 431 289
rect 433 285 437 289
rect 439 285 443 289
rect 445 285 449 289
rect 471 286 475 290
rect 489 286 493 290
rect 414 279 418 283
rect 420 279 424 283
rect 427 279 431 283
rect 433 279 437 283
rect 439 279 443 283
rect 445 279 449 283
rect 471 280 475 284
rect 489 280 493 284
rect 414 273 418 277
rect 420 273 424 277
rect 427 273 431 277
rect 433 273 437 277
rect 439 273 443 277
rect 445 273 449 277
rect 471 274 475 278
rect 489 274 493 278
rect 384 268 388 272
rect 397 268 401 272
rect 471 268 475 272
rect 489 268 493 272
rect 384 262 388 266
rect 397 262 401 266
rect 456 264 460 268
rect 471 262 475 266
rect 489 262 493 266
rect 456 254 460 258
rect 456 216 460 220
rect 384 208 388 212
rect 397 208 401 212
rect 456 206 460 210
rect 471 208 475 212
rect 489 208 493 212
rect 384 202 388 206
rect 397 202 401 206
rect 471 202 475 206
rect 489 202 493 206
rect 384 196 388 200
rect 397 196 401 200
rect 384 190 388 194
rect 397 190 401 194
rect 384 184 388 188
rect 397 184 401 188
rect 384 178 388 182
rect 397 178 401 182
rect 384 172 388 176
rect 397 172 401 176
rect 414 197 418 201
rect 420 197 424 201
rect 427 197 431 201
rect 433 197 437 201
rect 439 197 443 201
rect 445 197 449 201
rect 471 196 475 200
rect 489 196 493 200
rect 414 191 418 195
rect 420 191 424 195
rect 427 191 431 195
rect 433 191 437 195
rect 439 191 443 195
rect 445 191 449 195
rect 471 190 475 194
rect 489 190 493 194
rect 414 185 418 189
rect 420 185 424 189
rect 427 185 431 189
rect 433 185 437 189
rect 439 185 443 189
rect 445 185 449 189
rect 471 184 475 188
rect 489 184 493 188
rect 414 179 418 183
rect 420 179 424 183
rect 427 179 431 183
rect 433 179 437 183
rect 439 179 443 183
rect 445 179 449 183
rect 471 178 475 182
rect 489 178 493 182
rect 414 173 418 177
rect 420 173 424 177
rect 427 173 431 177
rect 433 173 437 177
rect 439 173 443 177
rect 445 173 449 177
rect 471 172 475 176
rect 489 172 493 176
<< electrodecap >>
rect 376 4143 408 4225
rect 381 4093 408 4143
rect 376 3965 408 4093
rect 381 3915 408 3965
rect 376 3669 408 3915
rect 381 3619 408 3669
rect 376 3491 408 3619
rect 381 3441 408 3491
rect 376 3195 408 3441
rect 381 3145 408 3195
rect 376 3017 408 3145
rect 381 2967 408 3017
rect 376 2721 408 2967
rect 381 2671 408 2721
rect 376 2543 408 2671
rect 381 2493 408 2543
rect 376 2247 408 2493
rect 381 2197 408 2247
rect 376 2069 408 2197
rect 381 2019 408 2069
rect 376 1773 408 2019
rect 381 1723 408 1773
rect 376 1595 408 1723
rect 381 1545 408 1595
rect 376 1299 408 1545
rect 381 1249 408 1299
rect 376 1121 408 1249
rect 381 1071 408 1121
rect 376 825 408 1071
rect 381 775 408 825
rect 376 647 408 775
rect 381 597 408 647
rect 376 351 408 597
rect 381 301 408 351
rect 376 173 408 301
rect 381 123 408 173
rect 376 41 408 123
rect 411 84 451 4182
rect 454 95 462 4171
rect 465 3965 501 4168
rect 465 3915 496 3965
rect 465 3669 501 3915
rect 465 3619 496 3669
rect 465 3491 501 3619
rect 465 3441 496 3491
rect 465 3195 501 3441
rect 465 3145 496 3195
rect 465 3017 501 3145
rect 465 2967 496 3017
rect 465 2721 501 2967
rect 465 2671 496 2721
rect 465 2543 501 2671
rect 465 2493 496 2543
rect 465 2247 501 2493
rect 465 2197 496 2247
rect 465 2069 501 2197
rect 465 2019 496 2069
rect 465 1773 501 2019
rect 465 1723 496 1773
rect 465 1595 501 1723
rect 465 1545 496 1595
rect 465 1299 501 1545
rect 465 1249 496 1299
rect 465 1121 501 1249
rect 465 1071 496 1121
rect 465 825 501 1071
rect 465 775 496 825
rect 465 647 501 775
rect 465 597 496 647
rect 465 351 501 597
rect 465 301 496 351
rect 465 98 501 301
<< psubstratepdiff >>
rect 364 4262 370 4263
rect 364 4258 365 4262
rect 369 4258 370 4262
rect 364 4256 370 4258
rect 364 4252 365 4256
rect 369 4252 370 4256
rect 364 4250 370 4252
rect 364 4246 365 4250
rect 369 4246 370 4250
rect 364 4244 370 4246
rect 364 4240 365 4244
rect 369 4240 370 4244
rect 364 4238 370 4240
rect 364 4234 365 4238
rect 369 4234 370 4238
rect 364 4232 370 4234
rect 364 4228 365 4232
rect 369 4228 370 4232
rect 364 4226 370 4228
rect 364 4222 365 4226
rect 369 4222 370 4226
rect 364 4220 370 4222
rect 364 4216 365 4220
rect 369 4216 370 4220
rect 364 4214 370 4216
rect 364 4210 365 4214
rect 369 4210 370 4214
rect 364 4208 370 4210
rect 364 4204 365 4208
rect 369 4204 370 4208
rect 364 4202 370 4204
rect 364 4198 365 4202
rect 369 4198 370 4202
rect 364 4196 370 4198
rect 364 4192 365 4196
rect 369 4192 370 4196
rect 364 4190 370 4192
rect 364 4186 365 4190
rect 369 4186 370 4190
rect 364 4184 370 4186
rect 364 4180 365 4184
rect 369 4180 370 4184
rect 364 4178 370 4180
rect 364 4174 365 4178
rect 369 4174 370 4178
rect 364 4172 370 4174
rect 364 4168 365 4172
rect 369 4168 370 4172
rect 364 4166 370 4168
rect 364 4162 365 4166
rect 369 4162 370 4166
rect 364 4160 370 4162
rect 364 4156 365 4160
rect 369 4156 370 4160
rect 364 4154 370 4156
rect 364 4150 365 4154
rect 369 4150 370 4154
rect 364 4148 370 4150
rect 364 4144 365 4148
rect 369 4144 370 4148
rect 364 4142 370 4144
rect 364 4138 365 4142
rect 369 4138 370 4142
rect 364 4136 370 4138
rect 364 4132 365 4136
rect 369 4132 370 4136
rect 364 4130 370 4132
rect 364 4126 365 4130
rect 369 4126 370 4130
rect 364 4124 370 4126
rect 364 4120 365 4124
rect 369 4120 370 4124
rect 364 4118 370 4120
rect 364 4114 365 4118
rect 369 4114 370 4118
rect 364 4112 370 4114
rect 364 4108 365 4112
rect 369 4108 370 4112
rect 364 4106 370 4108
rect 364 4102 365 4106
rect 369 4102 370 4106
rect 364 4100 370 4102
rect 364 4096 365 4100
rect 369 4096 370 4100
rect 364 4094 370 4096
rect 364 4090 365 4094
rect 369 4090 370 4094
rect 364 4088 370 4090
rect 364 4084 365 4088
rect 369 4084 370 4088
rect 364 4082 370 4084
rect 364 4078 365 4082
rect 369 4078 370 4082
rect 364 4076 370 4078
rect 364 4072 365 4076
rect 369 4072 370 4076
rect 364 4070 370 4072
rect 364 4066 365 4070
rect 369 4066 370 4070
rect 364 4064 370 4066
rect 364 4060 365 4064
rect 369 4060 370 4064
rect 364 4058 370 4060
rect 364 4054 365 4058
rect 369 4054 370 4058
rect 364 4052 370 4054
rect 364 4048 365 4052
rect 369 4048 370 4052
rect 364 4046 370 4048
rect 364 4042 365 4046
rect 369 4042 370 4046
rect 364 4016 370 4042
rect 364 4012 365 4016
rect 369 4012 370 4016
rect 364 4010 370 4012
rect 364 4006 365 4010
rect 369 4006 370 4010
rect 364 4004 370 4006
rect 364 4000 365 4004
rect 369 4000 370 4004
rect 364 3998 370 4000
rect 364 3994 365 3998
rect 369 3994 370 3998
rect 364 3992 370 3994
rect 364 3988 365 3992
rect 369 3988 370 3992
rect 364 3986 370 3988
rect 364 3982 365 3986
rect 369 3982 370 3986
rect 364 3980 370 3982
rect 364 3976 365 3980
rect 369 3976 370 3980
rect 364 3974 370 3976
rect 364 3970 365 3974
rect 369 3970 370 3974
rect 364 3968 370 3970
rect 364 3964 365 3968
rect 369 3964 370 3968
rect 364 3962 370 3964
rect 364 3958 365 3962
rect 369 3958 370 3962
rect 364 3956 370 3958
rect 364 3952 365 3956
rect 369 3952 370 3956
rect 364 3950 370 3952
rect 364 3946 365 3950
rect 369 3946 370 3950
rect 364 3944 370 3946
rect 364 3940 365 3944
rect 369 3940 370 3944
rect 364 3938 370 3940
rect 364 3934 365 3938
rect 369 3934 370 3938
rect 364 3932 370 3934
rect 364 3928 365 3932
rect 369 3928 370 3932
rect 364 3926 370 3928
rect 364 3922 365 3926
rect 369 3922 370 3926
rect 364 3920 370 3922
rect 364 3916 365 3920
rect 369 3916 370 3920
rect 364 3914 370 3916
rect 364 3910 365 3914
rect 369 3910 370 3914
rect 364 3908 370 3910
rect 364 3904 365 3908
rect 369 3904 370 3908
rect 364 3902 370 3904
rect 364 3898 365 3902
rect 369 3898 370 3902
rect 364 3896 370 3898
rect 364 3892 365 3896
rect 369 3892 370 3896
rect 364 3890 370 3892
rect 364 3886 365 3890
rect 369 3886 370 3890
rect 364 3884 370 3886
rect 364 3880 365 3884
rect 369 3880 370 3884
rect 364 3878 370 3880
rect 364 3874 365 3878
rect 369 3874 370 3878
rect 364 3872 370 3874
rect 364 3868 365 3872
rect 369 3868 370 3872
rect 364 3866 370 3868
rect 364 3862 365 3866
rect 369 3862 370 3866
rect 364 3860 370 3862
rect 364 3856 365 3860
rect 369 3856 370 3860
rect 364 3854 370 3856
rect 364 3850 365 3854
rect 369 3850 370 3854
rect 364 3848 370 3850
rect 364 3844 365 3848
rect 369 3844 370 3848
rect 364 3842 370 3844
rect 364 3838 365 3842
rect 369 3838 370 3842
rect 364 3836 370 3838
rect 364 3832 365 3836
rect 369 3832 370 3836
rect 364 3830 370 3832
rect 364 3826 365 3830
rect 369 3826 370 3830
rect 364 3824 370 3826
rect 364 3820 365 3824
rect 369 3820 370 3824
rect 364 3818 370 3820
rect 364 3814 365 3818
rect 369 3814 370 3818
rect 364 3812 370 3814
rect 364 3808 365 3812
rect 369 3808 370 3812
rect 364 3806 370 3808
rect 364 3802 365 3806
rect 369 3802 370 3806
rect 364 3800 370 3802
rect 364 3796 365 3800
rect 369 3796 370 3800
rect 364 3795 370 3796
rect 2 3794 370 3795
rect 2 3790 5 3794
rect 9 3790 11 3794
rect 15 3790 17 3794
rect 21 3790 23 3794
rect 27 3790 29 3794
rect 33 3790 35 3794
rect 39 3790 41 3794
rect 45 3790 47 3794
rect 51 3790 53 3794
rect 57 3790 59 3794
rect 63 3790 65 3794
rect 69 3790 71 3794
rect 75 3790 77 3794
rect 81 3790 83 3794
rect 87 3790 89 3794
rect 93 3790 95 3794
rect 99 3790 101 3794
rect 105 3790 107 3794
rect 111 3790 113 3794
rect 117 3790 119 3794
rect 123 3790 125 3794
rect 129 3790 131 3794
rect 135 3790 137 3794
rect 141 3790 143 3794
rect 147 3790 149 3794
rect 153 3790 155 3794
rect 159 3790 161 3794
rect 165 3790 167 3794
rect 171 3790 173 3794
rect 177 3790 179 3794
rect 183 3790 185 3794
rect 189 3790 191 3794
rect 195 3790 197 3794
rect 201 3790 203 3794
rect 207 3790 209 3794
rect 213 3790 215 3794
rect 219 3790 221 3794
rect 225 3790 227 3794
rect 231 3790 233 3794
rect 237 3790 239 3794
rect 243 3790 245 3794
rect 249 3790 251 3794
rect 255 3790 257 3794
rect 261 3790 263 3794
rect 267 3790 269 3794
rect 273 3790 275 3794
rect 279 3790 281 3794
rect 285 3790 287 3794
rect 291 3790 293 3794
rect 297 3790 299 3794
rect 303 3790 305 3794
rect 309 3790 311 3794
rect 315 3790 317 3794
rect 321 3790 323 3794
rect 327 3790 329 3794
rect 333 3790 335 3794
rect 339 3790 341 3794
rect 345 3790 347 3794
rect 351 3790 353 3794
rect 357 3790 359 3794
rect 363 3790 365 3794
rect 369 3790 370 3794
rect 2 3789 370 3790
rect 364 3788 370 3789
rect 364 3784 365 3788
rect 369 3784 370 3788
rect 364 3782 370 3784
rect 364 3778 365 3782
rect 369 3778 370 3782
rect 364 3776 370 3778
rect 364 3772 365 3776
rect 369 3772 370 3776
rect 364 3770 370 3772
rect 364 3766 365 3770
rect 369 3766 370 3770
rect 364 3764 370 3766
rect 364 3760 365 3764
rect 369 3760 370 3764
rect 364 3758 370 3760
rect 364 3754 365 3758
rect 369 3754 370 3758
rect 364 3752 370 3754
rect 364 3748 365 3752
rect 369 3748 370 3752
rect 364 3746 370 3748
rect 364 3742 365 3746
rect 369 3742 370 3746
rect 364 3740 370 3742
rect 364 3736 365 3740
rect 369 3736 370 3740
rect 364 3734 370 3736
rect 364 3730 365 3734
rect 369 3730 370 3734
rect 364 3728 370 3730
rect 364 3724 365 3728
rect 369 3724 370 3728
rect 364 3722 370 3724
rect 364 3718 365 3722
rect 369 3718 370 3722
rect 364 3716 370 3718
rect 364 3712 365 3716
rect 369 3712 370 3716
rect 364 3710 370 3712
rect 364 3706 365 3710
rect 369 3706 370 3710
rect 364 3704 370 3706
rect 364 3700 365 3704
rect 369 3700 370 3704
rect 364 3698 370 3700
rect 364 3694 365 3698
rect 369 3694 370 3698
rect 364 3692 370 3694
rect 364 3688 365 3692
rect 369 3688 370 3692
rect 364 3686 370 3688
rect 364 3682 365 3686
rect 369 3682 370 3686
rect 364 3680 370 3682
rect 364 3676 365 3680
rect 369 3676 370 3680
rect 364 3674 370 3676
rect 364 3670 365 3674
rect 369 3670 370 3674
rect 364 3668 370 3670
rect 364 3664 365 3668
rect 369 3664 370 3668
rect 364 3662 370 3664
rect 364 3658 365 3662
rect 369 3658 370 3662
rect 364 3656 370 3658
rect 364 3652 365 3656
rect 369 3652 370 3656
rect 364 3650 370 3652
rect 364 3646 365 3650
rect 369 3646 370 3650
rect 364 3644 370 3646
rect 364 3640 365 3644
rect 369 3640 370 3644
rect 364 3638 370 3640
rect 364 3634 365 3638
rect 369 3634 370 3638
rect 364 3632 370 3634
rect 364 3628 365 3632
rect 369 3628 370 3632
rect 364 3626 370 3628
rect 364 3622 365 3626
rect 369 3622 370 3626
rect 364 3620 370 3622
rect 364 3616 365 3620
rect 369 3616 370 3620
rect 364 3614 370 3616
rect 364 3610 365 3614
rect 369 3610 370 3614
rect 364 3608 370 3610
rect 364 3604 365 3608
rect 369 3604 370 3608
rect 364 3602 370 3604
rect 364 3598 365 3602
rect 369 3598 370 3602
rect 364 3596 370 3598
rect 364 3592 365 3596
rect 369 3592 370 3596
rect 364 3590 370 3592
rect 364 3586 365 3590
rect 369 3586 370 3590
rect 364 3584 370 3586
rect 364 3580 365 3584
rect 369 3580 370 3584
rect 364 3578 370 3580
rect 364 3574 365 3578
rect 369 3574 370 3578
rect 364 3572 370 3574
rect 364 3568 365 3572
rect 369 3568 370 3572
rect 364 3542 370 3568
rect 364 3538 365 3542
rect 369 3538 370 3542
rect 364 3536 370 3538
rect 364 3532 365 3536
rect 369 3532 370 3536
rect 364 3530 370 3532
rect 364 3526 365 3530
rect 369 3526 370 3530
rect 364 3524 370 3526
rect 364 3520 365 3524
rect 369 3520 370 3524
rect 364 3518 370 3520
rect 364 3514 365 3518
rect 369 3514 370 3518
rect 364 3512 370 3514
rect 364 3508 365 3512
rect 369 3508 370 3512
rect 364 3506 370 3508
rect 364 3502 365 3506
rect 369 3502 370 3506
rect 364 3500 370 3502
rect 364 3496 365 3500
rect 369 3496 370 3500
rect 364 3494 370 3496
rect 364 3490 365 3494
rect 369 3490 370 3494
rect 364 3488 370 3490
rect 364 3484 365 3488
rect 369 3484 370 3488
rect 364 3482 370 3484
rect 364 3478 365 3482
rect 369 3478 370 3482
rect 364 3476 370 3478
rect 364 3472 365 3476
rect 369 3472 370 3476
rect 364 3470 370 3472
rect 364 3466 365 3470
rect 369 3466 370 3470
rect 364 3464 370 3466
rect 364 3460 365 3464
rect 369 3460 370 3464
rect 364 3458 370 3460
rect 364 3454 365 3458
rect 369 3454 370 3458
rect 364 3452 370 3454
rect 364 3448 365 3452
rect 369 3448 370 3452
rect 364 3446 370 3448
rect 364 3442 365 3446
rect 369 3442 370 3446
rect 364 3440 370 3442
rect 364 3436 365 3440
rect 369 3436 370 3440
rect 364 3434 370 3436
rect 364 3430 365 3434
rect 369 3430 370 3434
rect 364 3428 370 3430
rect 364 3424 365 3428
rect 369 3424 370 3428
rect 364 3422 370 3424
rect 364 3418 365 3422
rect 369 3418 370 3422
rect 364 3416 370 3418
rect 364 3412 365 3416
rect 369 3412 370 3416
rect 364 3410 370 3412
rect 364 3406 365 3410
rect 369 3406 370 3410
rect 364 3404 370 3406
rect 364 3400 365 3404
rect 369 3400 370 3404
rect 364 3398 370 3400
rect 364 3394 365 3398
rect 369 3394 370 3398
rect 364 3392 370 3394
rect 364 3388 365 3392
rect 369 3388 370 3392
rect 364 3386 370 3388
rect 364 3382 365 3386
rect 369 3382 370 3386
rect 364 3380 370 3382
rect 364 3376 365 3380
rect 369 3376 370 3380
rect 364 3374 370 3376
rect 364 3370 365 3374
rect 369 3370 370 3374
rect 364 3368 370 3370
rect 364 3364 365 3368
rect 369 3364 370 3368
rect 364 3362 370 3364
rect 364 3358 365 3362
rect 369 3358 370 3362
rect 364 3356 370 3358
rect 364 3352 365 3356
rect 369 3352 370 3356
rect 364 3350 370 3352
rect 364 3346 365 3350
rect 369 3346 370 3350
rect 364 3344 370 3346
rect 364 3340 365 3344
rect 369 3340 370 3344
rect 364 3338 370 3340
rect 364 3334 365 3338
rect 369 3334 370 3338
rect 364 3332 370 3334
rect 364 3328 365 3332
rect 369 3328 370 3332
rect 364 3326 370 3328
rect 364 3322 365 3326
rect 369 3322 370 3326
rect 364 3321 370 3322
rect 2 3320 370 3321
rect 2 3316 5 3320
rect 9 3316 11 3320
rect 15 3316 17 3320
rect 21 3316 23 3320
rect 27 3316 29 3320
rect 33 3316 35 3320
rect 39 3316 41 3320
rect 45 3316 47 3320
rect 51 3316 53 3320
rect 57 3316 59 3320
rect 63 3316 65 3320
rect 69 3316 71 3320
rect 75 3316 77 3320
rect 81 3316 83 3320
rect 87 3316 89 3320
rect 93 3316 95 3320
rect 99 3316 101 3320
rect 105 3316 107 3320
rect 111 3316 113 3320
rect 117 3316 119 3320
rect 123 3316 125 3320
rect 129 3316 131 3320
rect 135 3316 137 3320
rect 141 3316 143 3320
rect 147 3316 149 3320
rect 153 3316 155 3320
rect 159 3316 161 3320
rect 165 3316 167 3320
rect 171 3316 173 3320
rect 177 3316 179 3320
rect 183 3316 185 3320
rect 189 3316 191 3320
rect 195 3316 197 3320
rect 201 3316 203 3320
rect 207 3316 209 3320
rect 213 3316 215 3320
rect 219 3316 221 3320
rect 225 3316 227 3320
rect 231 3316 233 3320
rect 237 3316 239 3320
rect 243 3316 245 3320
rect 249 3316 251 3320
rect 255 3316 257 3320
rect 261 3316 263 3320
rect 267 3316 269 3320
rect 273 3316 275 3320
rect 279 3316 281 3320
rect 285 3316 287 3320
rect 291 3316 293 3320
rect 297 3316 299 3320
rect 303 3316 305 3320
rect 309 3316 311 3320
rect 315 3316 317 3320
rect 321 3316 323 3320
rect 327 3316 329 3320
rect 333 3316 335 3320
rect 339 3316 341 3320
rect 345 3316 347 3320
rect 351 3316 353 3320
rect 357 3316 359 3320
rect 363 3316 365 3320
rect 369 3316 370 3320
rect 2 3315 370 3316
rect 364 3314 370 3315
rect 364 3310 365 3314
rect 369 3310 370 3314
rect 364 3308 370 3310
rect 364 3304 365 3308
rect 369 3304 370 3308
rect 364 3302 370 3304
rect 364 3298 365 3302
rect 369 3298 370 3302
rect 364 3296 370 3298
rect 364 3292 365 3296
rect 369 3292 370 3296
rect 364 3290 370 3292
rect 364 3286 365 3290
rect 369 3286 370 3290
rect 364 3284 370 3286
rect 364 3280 365 3284
rect 369 3280 370 3284
rect 364 3278 370 3280
rect 364 3274 365 3278
rect 369 3274 370 3278
rect 364 3272 370 3274
rect 364 3268 365 3272
rect 369 3268 370 3272
rect 364 3266 370 3268
rect 364 3262 365 3266
rect 369 3262 370 3266
rect 364 3260 370 3262
rect 364 3256 365 3260
rect 369 3256 370 3260
rect 364 3254 370 3256
rect 364 3250 365 3254
rect 369 3250 370 3254
rect 364 3248 370 3250
rect 364 3244 365 3248
rect 369 3244 370 3248
rect 364 3242 370 3244
rect 364 3238 365 3242
rect 369 3238 370 3242
rect 364 3236 370 3238
rect 364 3232 365 3236
rect 369 3232 370 3236
rect 364 3230 370 3232
rect 364 3226 365 3230
rect 369 3226 370 3230
rect 364 3224 370 3226
rect 364 3220 365 3224
rect 369 3220 370 3224
rect 364 3218 370 3220
rect 364 3214 365 3218
rect 369 3214 370 3218
rect 364 3212 370 3214
rect 364 3208 365 3212
rect 369 3208 370 3212
rect 364 3206 370 3208
rect 364 3202 365 3206
rect 369 3202 370 3206
rect 364 3200 370 3202
rect 364 3196 365 3200
rect 369 3196 370 3200
rect 364 3194 370 3196
rect 364 3190 365 3194
rect 369 3190 370 3194
rect 364 3188 370 3190
rect 364 3184 365 3188
rect 369 3184 370 3188
rect 364 3182 370 3184
rect 364 3178 365 3182
rect 369 3178 370 3182
rect 364 3176 370 3178
rect 364 3172 365 3176
rect 369 3172 370 3176
rect 364 3170 370 3172
rect 364 3166 365 3170
rect 369 3166 370 3170
rect 364 3164 370 3166
rect 364 3160 365 3164
rect 369 3160 370 3164
rect 364 3158 370 3160
rect 364 3154 365 3158
rect 369 3154 370 3158
rect 364 3152 370 3154
rect 364 3148 365 3152
rect 369 3148 370 3152
rect 364 3146 370 3148
rect 364 3142 365 3146
rect 369 3142 370 3146
rect 364 3140 370 3142
rect 364 3136 365 3140
rect 369 3136 370 3140
rect 364 3134 370 3136
rect 364 3130 365 3134
rect 369 3130 370 3134
rect 364 3128 370 3130
rect 364 3124 365 3128
rect 369 3124 370 3128
rect 364 3122 370 3124
rect 364 3118 365 3122
rect 369 3118 370 3122
rect 364 3116 370 3118
rect 364 3112 365 3116
rect 369 3112 370 3116
rect 364 3110 370 3112
rect 364 3106 365 3110
rect 369 3106 370 3110
rect 364 3104 370 3106
rect 364 3100 365 3104
rect 369 3100 370 3104
rect 364 3098 370 3100
rect 364 3094 365 3098
rect 369 3094 370 3098
rect 364 3068 370 3094
rect 364 3064 365 3068
rect 369 3064 370 3068
rect 364 3062 370 3064
rect 364 3058 365 3062
rect 369 3058 370 3062
rect 364 3056 370 3058
rect 364 3052 365 3056
rect 369 3052 370 3056
rect 364 3050 370 3052
rect 364 3046 365 3050
rect 369 3046 370 3050
rect 364 3044 370 3046
rect 364 3040 365 3044
rect 369 3040 370 3044
rect 364 3038 370 3040
rect 364 3034 365 3038
rect 369 3034 370 3038
rect 364 3032 370 3034
rect 364 3028 365 3032
rect 369 3028 370 3032
rect 364 3026 370 3028
rect 364 3022 365 3026
rect 369 3022 370 3026
rect 364 3020 370 3022
rect 364 3016 365 3020
rect 369 3016 370 3020
rect 364 3014 370 3016
rect 364 3010 365 3014
rect 369 3010 370 3014
rect 364 3008 370 3010
rect 364 3004 365 3008
rect 369 3004 370 3008
rect 364 3002 370 3004
rect 364 2998 365 3002
rect 369 2998 370 3002
rect 364 2996 370 2998
rect 364 2992 365 2996
rect 369 2992 370 2996
rect 364 2990 370 2992
rect 364 2986 365 2990
rect 369 2986 370 2990
rect 364 2984 370 2986
rect 364 2980 365 2984
rect 369 2980 370 2984
rect 364 2978 370 2980
rect 364 2974 365 2978
rect 369 2974 370 2978
rect 364 2972 370 2974
rect 364 2968 365 2972
rect 369 2968 370 2972
rect 364 2966 370 2968
rect 364 2962 365 2966
rect 369 2962 370 2966
rect 364 2960 370 2962
rect 364 2956 365 2960
rect 369 2956 370 2960
rect 364 2954 370 2956
rect 364 2950 365 2954
rect 369 2950 370 2954
rect 364 2948 370 2950
rect 364 2944 365 2948
rect 369 2944 370 2948
rect 364 2942 370 2944
rect 364 2938 365 2942
rect 369 2938 370 2942
rect 364 2936 370 2938
rect 364 2932 365 2936
rect 369 2932 370 2936
rect 364 2930 370 2932
rect 364 2926 365 2930
rect 369 2926 370 2930
rect 364 2924 370 2926
rect 364 2920 365 2924
rect 369 2920 370 2924
rect 364 2918 370 2920
rect 364 2914 365 2918
rect 369 2914 370 2918
rect 364 2912 370 2914
rect 364 2908 365 2912
rect 369 2908 370 2912
rect 364 2906 370 2908
rect 364 2902 365 2906
rect 369 2902 370 2906
rect 364 2900 370 2902
rect 364 2896 365 2900
rect 369 2896 370 2900
rect 364 2894 370 2896
rect 364 2890 365 2894
rect 369 2890 370 2894
rect 364 2888 370 2890
rect 364 2884 365 2888
rect 369 2884 370 2888
rect 364 2882 370 2884
rect 364 2878 365 2882
rect 369 2878 370 2882
rect 364 2876 370 2878
rect 364 2872 365 2876
rect 369 2872 370 2876
rect 364 2870 370 2872
rect 364 2866 365 2870
rect 369 2866 370 2870
rect 364 2864 370 2866
rect 364 2860 365 2864
rect 369 2860 370 2864
rect 364 2858 370 2860
rect 364 2854 365 2858
rect 369 2854 370 2858
rect 364 2852 370 2854
rect 364 2848 365 2852
rect 369 2848 370 2852
rect 364 2847 370 2848
rect 2 2846 370 2847
rect 2 2842 5 2846
rect 9 2842 11 2846
rect 15 2842 17 2846
rect 21 2842 23 2846
rect 27 2842 29 2846
rect 33 2842 35 2846
rect 39 2842 41 2846
rect 45 2842 47 2846
rect 51 2842 53 2846
rect 57 2842 59 2846
rect 63 2842 65 2846
rect 69 2842 71 2846
rect 75 2842 77 2846
rect 81 2842 83 2846
rect 87 2842 89 2846
rect 93 2842 95 2846
rect 99 2842 101 2846
rect 105 2842 107 2846
rect 111 2842 113 2846
rect 117 2842 119 2846
rect 123 2842 125 2846
rect 129 2842 131 2846
rect 135 2842 137 2846
rect 141 2842 143 2846
rect 147 2842 149 2846
rect 153 2842 155 2846
rect 159 2842 161 2846
rect 165 2842 167 2846
rect 171 2842 173 2846
rect 177 2842 179 2846
rect 183 2842 185 2846
rect 189 2842 191 2846
rect 195 2842 197 2846
rect 201 2842 203 2846
rect 207 2842 209 2846
rect 213 2842 215 2846
rect 219 2842 221 2846
rect 225 2842 227 2846
rect 231 2842 233 2846
rect 237 2842 239 2846
rect 243 2842 245 2846
rect 249 2842 251 2846
rect 255 2842 257 2846
rect 261 2842 263 2846
rect 267 2842 269 2846
rect 273 2842 275 2846
rect 279 2842 281 2846
rect 285 2842 287 2846
rect 291 2842 293 2846
rect 297 2842 299 2846
rect 303 2842 305 2846
rect 309 2842 311 2846
rect 315 2842 317 2846
rect 321 2842 323 2846
rect 327 2842 329 2846
rect 333 2842 335 2846
rect 339 2842 341 2846
rect 345 2842 347 2846
rect 351 2842 353 2846
rect 357 2842 359 2846
rect 363 2842 365 2846
rect 369 2842 370 2846
rect 2 2841 370 2842
rect 364 2840 370 2841
rect 364 2836 365 2840
rect 369 2836 370 2840
rect 364 2834 370 2836
rect 364 2830 365 2834
rect 369 2830 370 2834
rect 364 2828 370 2830
rect 364 2824 365 2828
rect 369 2824 370 2828
rect 364 2822 370 2824
rect 364 2818 365 2822
rect 369 2818 370 2822
rect 364 2816 370 2818
rect 364 2812 365 2816
rect 369 2812 370 2816
rect 364 2810 370 2812
rect 364 2806 365 2810
rect 369 2806 370 2810
rect 364 2804 370 2806
rect 364 2800 365 2804
rect 369 2800 370 2804
rect 364 2798 370 2800
rect 364 2794 365 2798
rect 369 2794 370 2798
rect 364 2792 370 2794
rect 364 2788 365 2792
rect 369 2788 370 2792
rect 364 2786 370 2788
rect 364 2782 365 2786
rect 369 2782 370 2786
rect 364 2780 370 2782
rect 364 2776 365 2780
rect 369 2776 370 2780
rect 364 2774 370 2776
rect 364 2770 365 2774
rect 369 2770 370 2774
rect 364 2768 370 2770
rect 364 2764 365 2768
rect 369 2764 370 2768
rect 364 2762 370 2764
rect 364 2758 365 2762
rect 369 2758 370 2762
rect 364 2756 370 2758
rect 364 2752 365 2756
rect 369 2752 370 2756
rect 364 2750 370 2752
rect 364 2746 365 2750
rect 369 2746 370 2750
rect 364 2744 370 2746
rect 364 2740 365 2744
rect 369 2740 370 2744
rect 364 2738 370 2740
rect 364 2734 365 2738
rect 369 2734 370 2738
rect 364 2732 370 2734
rect 364 2728 365 2732
rect 369 2728 370 2732
rect 364 2726 370 2728
rect 364 2722 365 2726
rect 369 2722 370 2726
rect 364 2720 370 2722
rect 364 2716 365 2720
rect 369 2716 370 2720
rect 364 2714 370 2716
rect 364 2710 365 2714
rect 369 2710 370 2714
rect 364 2708 370 2710
rect 364 2704 365 2708
rect 369 2704 370 2708
rect 364 2702 370 2704
rect 364 2698 365 2702
rect 369 2698 370 2702
rect 364 2696 370 2698
rect 364 2692 365 2696
rect 369 2692 370 2696
rect 364 2690 370 2692
rect 364 2686 365 2690
rect 369 2686 370 2690
rect 364 2684 370 2686
rect 364 2680 365 2684
rect 369 2680 370 2684
rect 364 2678 370 2680
rect 364 2674 365 2678
rect 369 2674 370 2678
rect 364 2672 370 2674
rect 364 2668 365 2672
rect 369 2668 370 2672
rect 364 2666 370 2668
rect 364 2662 365 2666
rect 369 2662 370 2666
rect 364 2660 370 2662
rect 364 2656 365 2660
rect 369 2656 370 2660
rect 364 2654 370 2656
rect 364 2650 365 2654
rect 369 2650 370 2654
rect 364 2648 370 2650
rect 364 2644 365 2648
rect 369 2644 370 2648
rect 364 2642 370 2644
rect 364 2638 365 2642
rect 369 2638 370 2642
rect 364 2636 370 2638
rect 364 2632 365 2636
rect 369 2632 370 2636
rect 364 2630 370 2632
rect 364 2626 365 2630
rect 369 2626 370 2630
rect 364 2624 370 2626
rect 364 2620 365 2624
rect 369 2620 370 2624
rect 364 2594 370 2620
rect 364 2590 365 2594
rect 369 2590 370 2594
rect 364 2588 370 2590
rect 364 2584 365 2588
rect 369 2584 370 2588
rect 364 2582 370 2584
rect 364 2578 365 2582
rect 369 2578 370 2582
rect 364 2576 370 2578
rect 364 2572 365 2576
rect 369 2572 370 2576
rect 364 2570 370 2572
rect 364 2566 365 2570
rect 369 2566 370 2570
rect 364 2564 370 2566
rect 364 2560 365 2564
rect 369 2560 370 2564
rect 364 2558 370 2560
rect 364 2554 365 2558
rect 369 2554 370 2558
rect 364 2552 370 2554
rect 364 2548 365 2552
rect 369 2548 370 2552
rect 364 2546 370 2548
rect 364 2542 365 2546
rect 369 2542 370 2546
rect 364 2540 370 2542
rect 364 2536 365 2540
rect 369 2536 370 2540
rect 364 2534 370 2536
rect 364 2530 365 2534
rect 369 2530 370 2534
rect 364 2528 370 2530
rect 364 2524 365 2528
rect 369 2524 370 2528
rect 364 2522 370 2524
rect 364 2518 365 2522
rect 369 2518 370 2522
rect 364 2516 370 2518
rect 364 2512 365 2516
rect 369 2512 370 2516
rect 364 2510 370 2512
rect 364 2506 365 2510
rect 369 2506 370 2510
rect 364 2504 370 2506
rect 364 2500 365 2504
rect 369 2500 370 2504
rect 364 2498 370 2500
rect 364 2494 365 2498
rect 369 2494 370 2498
rect 364 2492 370 2494
rect 364 2488 365 2492
rect 369 2488 370 2492
rect 364 2486 370 2488
rect 364 2482 365 2486
rect 369 2482 370 2486
rect 364 2480 370 2482
rect 364 2476 365 2480
rect 369 2476 370 2480
rect 364 2474 370 2476
rect 364 2470 365 2474
rect 369 2470 370 2474
rect 364 2468 370 2470
rect 364 2464 365 2468
rect 369 2464 370 2468
rect 364 2462 370 2464
rect 364 2458 365 2462
rect 369 2458 370 2462
rect 364 2456 370 2458
rect 364 2452 365 2456
rect 369 2452 370 2456
rect 364 2450 370 2452
rect 364 2446 365 2450
rect 369 2446 370 2450
rect 364 2444 370 2446
rect 364 2440 365 2444
rect 369 2440 370 2444
rect 364 2438 370 2440
rect 364 2434 365 2438
rect 369 2434 370 2438
rect 364 2432 370 2434
rect 364 2428 365 2432
rect 369 2428 370 2432
rect 364 2426 370 2428
rect 364 2422 365 2426
rect 369 2422 370 2426
rect 364 2420 370 2422
rect 364 2416 365 2420
rect 369 2416 370 2420
rect 364 2414 370 2416
rect 364 2410 365 2414
rect 369 2410 370 2414
rect 364 2408 370 2410
rect 364 2404 365 2408
rect 369 2404 370 2408
rect 364 2402 370 2404
rect 364 2398 365 2402
rect 369 2398 370 2402
rect 364 2396 370 2398
rect 364 2392 365 2396
rect 369 2392 370 2396
rect 364 2390 370 2392
rect 364 2386 365 2390
rect 369 2386 370 2390
rect 364 2384 370 2386
rect 364 2380 365 2384
rect 369 2380 370 2384
rect 364 2378 370 2380
rect 364 2374 365 2378
rect 369 2374 370 2378
rect 364 2373 370 2374
rect 2 2372 370 2373
rect 2 2368 5 2372
rect 9 2368 11 2372
rect 15 2368 17 2372
rect 21 2368 23 2372
rect 27 2368 29 2372
rect 33 2368 35 2372
rect 39 2368 41 2372
rect 45 2368 47 2372
rect 51 2368 53 2372
rect 57 2368 59 2372
rect 63 2368 65 2372
rect 69 2368 71 2372
rect 75 2368 77 2372
rect 81 2368 83 2372
rect 87 2368 89 2372
rect 93 2368 95 2372
rect 99 2368 101 2372
rect 105 2368 107 2372
rect 111 2368 113 2372
rect 117 2368 119 2372
rect 123 2368 125 2372
rect 129 2368 131 2372
rect 135 2368 137 2372
rect 141 2368 143 2372
rect 147 2368 149 2372
rect 153 2368 155 2372
rect 159 2368 161 2372
rect 165 2368 167 2372
rect 171 2368 173 2372
rect 177 2368 179 2372
rect 183 2368 185 2372
rect 189 2368 191 2372
rect 195 2368 197 2372
rect 201 2368 203 2372
rect 207 2368 209 2372
rect 213 2368 215 2372
rect 219 2368 221 2372
rect 225 2368 227 2372
rect 231 2368 233 2372
rect 237 2368 239 2372
rect 243 2368 245 2372
rect 249 2368 251 2372
rect 255 2368 257 2372
rect 261 2368 263 2372
rect 267 2368 269 2372
rect 273 2368 275 2372
rect 279 2368 281 2372
rect 285 2368 287 2372
rect 291 2368 293 2372
rect 297 2368 299 2372
rect 303 2368 305 2372
rect 309 2368 311 2372
rect 315 2368 317 2372
rect 321 2368 323 2372
rect 327 2368 329 2372
rect 333 2368 335 2372
rect 339 2368 341 2372
rect 345 2368 347 2372
rect 351 2368 353 2372
rect 357 2368 359 2372
rect 363 2368 365 2372
rect 369 2368 370 2372
rect 2 2367 370 2368
rect 364 2366 370 2367
rect 364 2362 365 2366
rect 369 2362 370 2366
rect 364 2360 370 2362
rect 364 2356 365 2360
rect 369 2356 370 2360
rect 364 2354 370 2356
rect 364 2350 365 2354
rect 369 2350 370 2354
rect 364 2348 370 2350
rect 364 2344 365 2348
rect 369 2344 370 2348
rect 364 2342 370 2344
rect 364 2338 365 2342
rect 369 2338 370 2342
rect 364 2336 370 2338
rect 364 2332 365 2336
rect 369 2332 370 2336
rect 364 2330 370 2332
rect 364 2326 365 2330
rect 369 2326 370 2330
rect 364 2324 370 2326
rect 364 2320 365 2324
rect 369 2320 370 2324
rect 364 2318 370 2320
rect 364 2314 365 2318
rect 369 2314 370 2318
rect 364 2312 370 2314
rect 364 2308 365 2312
rect 369 2308 370 2312
rect 364 2306 370 2308
rect 364 2302 365 2306
rect 369 2302 370 2306
rect 364 2300 370 2302
rect 364 2296 365 2300
rect 369 2296 370 2300
rect 364 2294 370 2296
rect 364 2290 365 2294
rect 369 2290 370 2294
rect 364 2288 370 2290
rect 364 2284 365 2288
rect 369 2284 370 2288
rect 364 2282 370 2284
rect 364 2278 365 2282
rect 369 2278 370 2282
rect 364 2276 370 2278
rect 364 2272 365 2276
rect 369 2272 370 2276
rect 364 2270 370 2272
rect 364 2266 365 2270
rect 369 2266 370 2270
rect 364 2264 370 2266
rect 364 2260 365 2264
rect 369 2260 370 2264
rect 364 2258 370 2260
rect 364 2254 365 2258
rect 369 2254 370 2258
rect 364 2252 370 2254
rect 364 2248 365 2252
rect 369 2248 370 2252
rect 364 2246 370 2248
rect 364 2242 365 2246
rect 369 2242 370 2246
rect 364 2240 370 2242
rect 364 2236 365 2240
rect 369 2236 370 2240
rect 364 2234 370 2236
rect 364 2230 365 2234
rect 369 2230 370 2234
rect 364 2228 370 2230
rect 364 2224 365 2228
rect 369 2224 370 2228
rect 364 2222 370 2224
rect 364 2218 365 2222
rect 369 2218 370 2222
rect 364 2216 370 2218
rect 364 2212 365 2216
rect 369 2212 370 2216
rect 364 2210 370 2212
rect 364 2206 365 2210
rect 369 2206 370 2210
rect 364 2204 370 2206
rect 364 2200 365 2204
rect 369 2200 370 2204
rect 364 2198 370 2200
rect 364 2194 365 2198
rect 369 2194 370 2198
rect 364 2192 370 2194
rect 364 2188 365 2192
rect 369 2188 370 2192
rect 364 2186 370 2188
rect 364 2182 365 2186
rect 369 2182 370 2186
rect 364 2180 370 2182
rect 364 2176 365 2180
rect 369 2176 370 2180
rect 364 2174 370 2176
rect 364 2170 365 2174
rect 369 2170 370 2174
rect 364 2168 370 2170
rect 364 2164 365 2168
rect 369 2164 370 2168
rect 364 2162 370 2164
rect 364 2158 365 2162
rect 369 2158 370 2162
rect 364 2156 370 2158
rect 364 2152 365 2156
rect 369 2152 370 2156
rect 364 2150 370 2152
rect 364 2146 365 2150
rect 369 2146 370 2150
rect 364 2120 370 2146
rect 364 2116 365 2120
rect 369 2116 370 2120
rect 364 2114 370 2116
rect 364 2110 365 2114
rect 369 2110 370 2114
rect 364 2108 370 2110
rect 364 2104 365 2108
rect 369 2104 370 2108
rect 364 2102 370 2104
rect 364 2098 365 2102
rect 369 2098 370 2102
rect 364 2096 370 2098
rect 364 2092 365 2096
rect 369 2092 370 2096
rect 364 2090 370 2092
rect 364 2086 365 2090
rect 369 2086 370 2090
rect 364 2084 370 2086
rect 364 2080 365 2084
rect 369 2080 370 2084
rect 364 2078 370 2080
rect 364 2074 365 2078
rect 369 2074 370 2078
rect 364 2072 370 2074
rect 364 2068 365 2072
rect 369 2068 370 2072
rect 364 2066 370 2068
rect 364 2062 365 2066
rect 369 2062 370 2066
rect 364 2060 370 2062
rect 364 2056 365 2060
rect 369 2056 370 2060
rect 364 2054 370 2056
rect 364 2050 365 2054
rect 369 2050 370 2054
rect 364 2048 370 2050
rect 364 2044 365 2048
rect 369 2044 370 2048
rect 364 2042 370 2044
rect 364 2038 365 2042
rect 369 2038 370 2042
rect 364 2036 370 2038
rect 364 2032 365 2036
rect 369 2032 370 2036
rect 364 2030 370 2032
rect 364 2026 365 2030
rect 369 2026 370 2030
rect 364 2024 370 2026
rect 364 2020 365 2024
rect 369 2020 370 2024
rect 364 2018 370 2020
rect 364 2014 365 2018
rect 369 2014 370 2018
rect 364 2012 370 2014
rect 364 2008 365 2012
rect 369 2008 370 2012
rect 364 2006 370 2008
rect 364 2002 365 2006
rect 369 2002 370 2006
rect 364 2000 370 2002
rect 364 1996 365 2000
rect 369 1996 370 2000
rect 364 1994 370 1996
rect 364 1990 365 1994
rect 369 1990 370 1994
rect 364 1988 370 1990
rect 364 1984 365 1988
rect 369 1984 370 1988
rect 364 1982 370 1984
rect 364 1978 365 1982
rect 369 1978 370 1982
rect 364 1976 370 1978
rect 364 1972 365 1976
rect 369 1972 370 1976
rect 364 1970 370 1972
rect 364 1966 365 1970
rect 369 1966 370 1970
rect 364 1964 370 1966
rect 364 1960 365 1964
rect 369 1960 370 1964
rect 364 1958 370 1960
rect 364 1954 365 1958
rect 369 1954 370 1958
rect 364 1952 370 1954
rect 364 1948 365 1952
rect 369 1948 370 1952
rect 364 1946 370 1948
rect 364 1942 365 1946
rect 369 1942 370 1946
rect 364 1940 370 1942
rect 364 1936 365 1940
rect 369 1936 370 1940
rect 364 1934 370 1936
rect 364 1930 365 1934
rect 369 1930 370 1934
rect 364 1928 370 1930
rect 364 1924 365 1928
rect 369 1924 370 1928
rect 364 1922 370 1924
rect 364 1918 365 1922
rect 369 1918 370 1922
rect 364 1916 370 1918
rect 364 1912 365 1916
rect 369 1912 370 1916
rect 364 1910 370 1912
rect 364 1906 365 1910
rect 369 1906 370 1910
rect 364 1904 370 1906
rect 364 1900 365 1904
rect 369 1900 370 1904
rect 364 1899 370 1900
rect 2 1898 370 1899
rect 2 1894 5 1898
rect 9 1894 11 1898
rect 15 1894 17 1898
rect 21 1894 23 1898
rect 27 1894 29 1898
rect 33 1894 35 1898
rect 39 1894 41 1898
rect 45 1894 47 1898
rect 51 1894 53 1898
rect 57 1894 59 1898
rect 63 1894 65 1898
rect 69 1894 71 1898
rect 75 1894 77 1898
rect 81 1894 83 1898
rect 87 1894 89 1898
rect 93 1894 95 1898
rect 99 1894 101 1898
rect 105 1894 107 1898
rect 111 1894 113 1898
rect 117 1894 119 1898
rect 123 1894 125 1898
rect 129 1894 131 1898
rect 135 1894 137 1898
rect 141 1894 143 1898
rect 147 1894 149 1898
rect 153 1894 155 1898
rect 159 1894 161 1898
rect 165 1894 167 1898
rect 171 1894 173 1898
rect 177 1894 179 1898
rect 183 1894 185 1898
rect 189 1894 191 1898
rect 195 1894 197 1898
rect 201 1894 203 1898
rect 207 1894 209 1898
rect 213 1894 215 1898
rect 219 1894 221 1898
rect 225 1894 227 1898
rect 231 1894 233 1898
rect 237 1894 239 1898
rect 243 1894 245 1898
rect 249 1894 251 1898
rect 255 1894 257 1898
rect 261 1894 263 1898
rect 267 1894 269 1898
rect 273 1894 275 1898
rect 279 1894 281 1898
rect 285 1894 287 1898
rect 291 1894 293 1898
rect 297 1894 299 1898
rect 303 1894 305 1898
rect 309 1894 311 1898
rect 315 1894 317 1898
rect 321 1894 323 1898
rect 327 1894 329 1898
rect 333 1894 335 1898
rect 339 1894 341 1898
rect 345 1894 347 1898
rect 351 1894 353 1898
rect 357 1894 359 1898
rect 363 1894 365 1898
rect 369 1894 370 1898
rect 2 1893 370 1894
rect 364 1892 370 1893
rect 364 1888 365 1892
rect 369 1888 370 1892
rect 364 1886 370 1888
rect 364 1882 365 1886
rect 369 1882 370 1886
rect 364 1880 370 1882
rect 364 1876 365 1880
rect 369 1876 370 1880
rect 364 1874 370 1876
rect 364 1870 365 1874
rect 369 1870 370 1874
rect 364 1868 370 1870
rect 364 1864 365 1868
rect 369 1864 370 1868
rect 364 1862 370 1864
rect 364 1858 365 1862
rect 369 1858 370 1862
rect 364 1856 370 1858
rect 364 1852 365 1856
rect 369 1852 370 1856
rect 364 1850 370 1852
rect 364 1846 365 1850
rect 369 1846 370 1850
rect 364 1844 370 1846
rect 364 1840 365 1844
rect 369 1840 370 1844
rect 364 1838 370 1840
rect 364 1834 365 1838
rect 369 1834 370 1838
rect 364 1832 370 1834
rect 364 1828 365 1832
rect 369 1828 370 1832
rect 364 1826 370 1828
rect 364 1822 365 1826
rect 369 1822 370 1826
rect 364 1820 370 1822
rect 364 1816 365 1820
rect 369 1816 370 1820
rect 364 1814 370 1816
rect 364 1810 365 1814
rect 369 1810 370 1814
rect 364 1808 370 1810
rect 364 1804 365 1808
rect 369 1804 370 1808
rect 364 1802 370 1804
rect 364 1798 365 1802
rect 369 1798 370 1802
rect 364 1796 370 1798
rect 364 1792 365 1796
rect 369 1792 370 1796
rect 364 1790 370 1792
rect 364 1786 365 1790
rect 369 1786 370 1790
rect 364 1784 370 1786
rect 364 1780 365 1784
rect 369 1780 370 1784
rect 364 1778 370 1780
rect 364 1774 365 1778
rect 369 1774 370 1778
rect 364 1772 370 1774
rect 364 1768 365 1772
rect 369 1768 370 1772
rect 364 1766 370 1768
rect 364 1762 365 1766
rect 369 1762 370 1766
rect 364 1760 370 1762
rect 364 1756 365 1760
rect 369 1756 370 1760
rect 364 1754 370 1756
rect 364 1750 365 1754
rect 369 1750 370 1754
rect 364 1748 370 1750
rect 364 1744 365 1748
rect 369 1744 370 1748
rect 364 1742 370 1744
rect 364 1738 365 1742
rect 369 1738 370 1742
rect 364 1736 370 1738
rect 364 1732 365 1736
rect 369 1732 370 1736
rect 364 1730 370 1732
rect 364 1726 365 1730
rect 369 1726 370 1730
rect 364 1724 370 1726
rect 364 1720 365 1724
rect 369 1720 370 1724
rect 364 1718 370 1720
rect 364 1714 365 1718
rect 369 1714 370 1718
rect 364 1712 370 1714
rect 364 1708 365 1712
rect 369 1708 370 1712
rect 364 1706 370 1708
rect 364 1702 365 1706
rect 369 1702 370 1706
rect 364 1700 370 1702
rect 364 1696 365 1700
rect 369 1696 370 1700
rect 364 1694 370 1696
rect 364 1690 365 1694
rect 369 1690 370 1694
rect 364 1688 370 1690
rect 364 1684 365 1688
rect 369 1684 370 1688
rect 364 1682 370 1684
rect 364 1678 365 1682
rect 369 1678 370 1682
rect 364 1676 370 1678
rect 364 1672 365 1676
rect 369 1672 370 1676
rect 364 1646 370 1672
rect 364 1642 365 1646
rect 369 1642 370 1646
rect 364 1640 370 1642
rect 364 1636 365 1640
rect 369 1636 370 1640
rect 364 1634 370 1636
rect 364 1630 365 1634
rect 369 1630 370 1634
rect 364 1628 370 1630
rect 364 1624 365 1628
rect 369 1624 370 1628
rect 364 1622 370 1624
rect 364 1618 365 1622
rect 369 1618 370 1622
rect 364 1616 370 1618
rect 364 1612 365 1616
rect 369 1612 370 1616
rect 364 1610 370 1612
rect 364 1606 365 1610
rect 369 1606 370 1610
rect 364 1604 370 1606
rect 364 1600 365 1604
rect 369 1600 370 1604
rect 364 1598 370 1600
rect 364 1594 365 1598
rect 369 1594 370 1598
rect 364 1592 370 1594
rect 364 1588 365 1592
rect 369 1588 370 1592
rect 364 1586 370 1588
rect 364 1582 365 1586
rect 369 1582 370 1586
rect 364 1580 370 1582
rect 364 1576 365 1580
rect 369 1576 370 1580
rect 364 1574 370 1576
rect 364 1570 365 1574
rect 369 1570 370 1574
rect 364 1568 370 1570
rect 364 1564 365 1568
rect 369 1564 370 1568
rect 364 1562 370 1564
rect 364 1558 365 1562
rect 369 1558 370 1562
rect 364 1556 370 1558
rect 364 1552 365 1556
rect 369 1552 370 1556
rect 364 1550 370 1552
rect 364 1546 365 1550
rect 369 1546 370 1550
rect 364 1544 370 1546
rect 364 1540 365 1544
rect 369 1540 370 1544
rect 364 1538 370 1540
rect 364 1534 365 1538
rect 369 1534 370 1538
rect 364 1532 370 1534
rect 364 1528 365 1532
rect 369 1528 370 1532
rect 364 1526 370 1528
rect 364 1522 365 1526
rect 369 1522 370 1526
rect 364 1520 370 1522
rect 364 1516 365 1520
rect 369 1516 370 1520
rect 364 1514 370 1516
rect 364 1510 365 1514
rect 369 1510 370 1514
rect 364 1508 370 1510
rect 364 1504 365 1508
rect 369 1504 370 1508
rect 364 1502 370 1504
rect 364 1498 365 1502
rect 369 1498 370 1502
rect 364 1496 370 1498
rect 364 1492 365 1496
rect 369 1492 370 1496
rect 364 1490 370 1492
rect 364 1486 365 1490
rect 369 1486 370 1490
rect 364 1484 370 1486
rect 364 1480 365 1484
rect 369 1480 370 1484
rect 364 1478 370 1480
rect 364 1474 365 1478
rect 369 1474 370 1478
rect 364 1472 370 1474
rect 364 1468 365 1472
rect 369 1468 370 1472
rect 364 1466 370 1468
rect 364 1462 365 1466
rect 369 1462 370 1466
rect 364 1460 370 1462
rect 364 1456 365 1460
rect 369 1456 370 1460
rect 364 1454 370 1456
rect 364 1450 365 1454
rect 369 1450 370 1454
rect 364 1448 370 1450
rect 364 1444 365 1448
rect 369 1444 370 1448
rect 364 1442 370 1444
rect 364 1438 365 1442
rect 369 1438 370 1442
rect 364 1436 370 1438
rect 364 1432 365 1436
rect 369 1432 370 1436
rect 364 1430 370 1432
rect 364 1426 365 1430
rect 369 1426 370 1430
rect 364 1425 370 1426
rect 2 1424 370 1425
rect 2 1420 5 1424
rect 9 1420 11 1424
rect 15 1420 17 1424
rect 21 1420 23 1424
rect 27 1420 29 1424
rect 33 1420 35 1424
rect 39 1420 41 1424
rect 45 1420 47 1424
rect 51 1420 53 1424
rect 57 1420 59 1424
rect 63 1420 65 1424
rect 69 1420 71 1424
rect 75 1420 77 1424
rect 81 1420 83 1424
rect 87 1420 89 1424
rect 93 1420 95 1424
rect 99 1420 101 1424
rect 105 1420 107 1424
rect 111 1420 113 1424
rect 117 1420 119 1424
rect 123 1420 125 1424
rect 129 1420 131 1424
rect 135 1420 137 1424
rect 141 1420 143 1424
rect 147 1420 149 1424
rect 153 1420 155 1424
rect 159 1420 161 1424
rect 165 1420 167 1424
rect 171 1420 173 1424
rect 177 1420 179 1424
rect 183 1420 185 1424
rect 189 1420 191 1424
rect 195 1420 197 1424
rect 201 1420 203 1424
rect 207 1420 209 1424
rect 213 1420 215 1424
rect 219 1420 221 1424
rect 225 1420 227 1424
rect 231 1420 233 1424
rect 237 1420 239 1424
rect 243 1420 245 1424
rect 249 1420 251 1424
rect 255 1420 257 1424
rect 261 1420 263 1424
rect 267 1420 269 1424
rect 273 1420 275 1424
rect 279 1420 281 1424
rect 285 1420 287 1424
rect 291 1420 293 1424
rect 297 1420 299 1424
rect 303 1420 305 1424
rect 309 1420 311 1424
rect 315 1420 317 1424
rect 321 1420 323 1424
rect 327 1420 329 1424
rect 333 1420 335 1424
rect 339 1420 341 1424
rect 345 1420 347 1424
rect 351 1420 353 1424
rect 357 1420 359 1424
rect 363 1420 365 1424
rect 369 1420 370 1424
rect 2 1419 370 1420
rect 364 1418 370 1419
rect 364 1414 365 1418
rect 369 1414 370 1418
rect 364 1412 370 1414
rect 364 1408 365 1412
rect 369 1408 370 1412
rect 364 1406 370 1408
rect 364 1402 365 1406
rect 369 1402 370 1406
rect 364 1400 370 1402
rect 364 1396 365 1400
rect 369 1396 370 1400
rect 364 1394 370 1396
rect 364 1390 365 1394
rect 369 1390 370 1394
rect 364 1388 370 1390
rect 364 1384 365 1388
rect 369 1384 370 1388
rect 364 1382 370 1384
rect 364 1378 365 1382
rect 369 1378 370 1382
rect 364 1376 370 1378
rect 364 1372 365 1376
rect 369 1372 370 1376
rect 364 1370 370 1372
rect 364 1366 365 1370
rect 369 1366 370 1370
rect 364 1364 370 1366
rect 364 1360 365 1364
rect 369 1360 370 1364
rect 364 1358 370 1360
rect 364 1354 365 1358
rect 369 1354 370 1358
rect 364 1352 370 1354
rect 364 1348 365 1352
rect 369 1348 370 1352
rect 364 1346 370 1348
rect 364 1342 365 1346
rect 369 1342 370 1346
rect 364 1340 370 1342
rect 364 1336 365 1340
rect 369 1336 370 1340
rect 364 1334 370 1336
rect 364 1330 365 1334
rect 369 1330 370 1334
rect 364 1328 370 1330
rect 364 1324 365 1328
rect 369 1324 370 1328
rect 364 1322 370 1324
rect 364 1318 365 1322
rect 369 1318 370 1322
rect 364 1316 370 1318
rect 364 1312 365 1316
rect 369 1312 370 1316
rect 364 1310 370 1312
rect 364 1306 365 1310
rect 369 1306 370 1310
rect 364 1304 370 1306
rect 364 1300 365 1304
rect 369 1300 370 1304
rect 364 1298 370 1300
rect 364 1294 365 1298
rect 369 1294 370 1298
rect 364 1292 370 1294
rect 364 1288 365 1292
rect 369 1288 370 1292
rect 364 1286 370 1288
rect 364 1282 365 1286
rect 369 1282 370 1286
rect 364 1280 370 1282
rect 364 1276 365 1280
rect 369 1276 370 1280
rect 364 1274 370 1276
rect 364 1270 365 1274
rect 369 1270 370 1274
rect 364 1268 370 1270
rect 364 1264 365 1268
rect 369 1264 370 1268
rect 364 1262 370 1264
rect 364 1258 365 1262
rect 369 1258 370 1262
rect 364 1256 370 1258
rect 364 1252 365 1256
rect 369 1252 370 1256
rect 364 1250 370 1252
rect 364 1246 365 1250
rect 369 1246 370 1250
rect 364 1244 370 1246
rect 364 1240 365 1244
rect 369 1240 370 1244
rect 364 1238 370 1240
rect 364 1234 365 1238
rect 369 1234 370 1238
rect 364 1232 370 1234
rect 364 1228 365 1232
rect 369 1228 370 1232
rect 364 1226 370 1228
rect 364 1222 365 1226
rect 369 1222 370 1226
rect 364 1220 370 1222
rect 364 1216 365 1220
rect 369 1216 370 1220
rect 364 1214 370 1216
rect 364 1210 365 1214
rect 369 1210 370 1214
rect 364 1208 370 1210
rect 364 1204 365 1208
rect 369 1204 370 1208
rect 364 1202 370 1204
rect 364 1198 365 1202
rect 369 1198 370 1202
rect 364 1172 370 1198
rect 364 1168 365 1172
rect 369 1168 370 1172
rect 364 1166 370 1168
rect 364 1162 365 1166
rect 369 1162 370 1166
rect 364 1160 370 1162
rect 364 1156 365 1160
rect 369 1156 370 1160
rect 364 1154 370 1156
rect 364 1150 365 1154
rect 369 1150 370 1154
rect 364 1148 370 1150
rect 364 1144 365 1148
rect 369 1144 370 1148
rect 364 1142 370 1144
rect 364 1138 365 1142
rect 369 1138 370 1142
rect 364 1136 370 1138
rect 364 1132 365 1136
rect 369 1132 370 1136
rect 364 1130 370 1132
rect 364 1126 365 1130
rect 369 1126 370 1130
rect 364 1124 370 1126
rect 364 1120 365 1124
rect 369 1120 370 1124
rect 364 1118 370 1120
rect 364 1114 365 1118
rect 369 1114 370 1118
rect 364 1112 370 1114
rect 364 1108 365 1112
rect 369 1108 370 1112
rect 364 1106 370 1108
rect 364 1102 365 1106
rect 369 1102 370 1106
rect 364 1100 370 1102
rect 364 1096 365 1100
rect 369 1096 370 1100
rect 364 1094 370 1096
rect 364 1090 365 1094
rect 369 1090 370 1094
rect 364 1088 370 1090
rect 364 1084 365 1088
rect 369 1084 370 1088
rect 364 1082 370 1084
rect 364 1078 365 1082
rect 369 1078 370 1082
rect 364 1076 370 1078
rect 364 1072 365 1076
rect 369 1072 370 1076
rect 364 1070 370 1072
rect 364 1066 365 1070
rect 369 1066 370 1070
rect 364 1064 370 1066
rect 364 1060 365 1064
rect 369 1060 370 1064
rect 364 1058 370 1060
rect 364 1054 365 1058
rect 369 1054 370 1058
rect 364 1052 370 1054
rect 364 1048 365 1052
rect 369 1048 370 1052
rect 364 1046 370 1048
rect 364 1042 365 1046
rect 369 1042 370 1046
rect 364 1040 370 1042
rect 364 1036 365 1040
rect 369 1036 370 1040
rect 364 1034 370 1036
rect 364 1030 365 1034
rect 369 1030 370 1034
rect 364 1028 370 1030
rect 364 1024 365 1028
rect 369 1024 370 1028
rect 364 1022 370 1024
rect 364 1018 365 1022
rect 369 1018 370 1022
rect 364 1016 370 1018
rect 364 1012 365 1016
rect 369 1012 370 1016
rect 364 1010 370 1012
rect 364 1006 365 1010
rect 369 1006 370 1010
rect 364 1004 370 1006
rect 364 1000 365 1004
rect 369 1000 370 1004
rect 364 998 370 1000
rect 364 994 365 998
rect 369 994 370 998
rect 364 992 370 994
rect 364 988 365 992
rect 369 988 370 992
rect 364 986 370 988
rect 364 982 365 986
rect 369 982 370 986
rect 364 980 370 982
rect 364 976 365 980
rect 369 976 370 980
rect 364 974 370 976
rect 364 970 365 974
rect 369 970 370 974
rect 364 968 370 970
rect 364 964 365 968
rect 369 964 370 968
rect 364 962 370 964
rect 364 958 365 962
rect 369 958 370 962
rect 364 956 370 958
rect 364 952 365 956
rect 369 952 370 956
rect 364 951 370 952
rect 2 950 370 951
rect 2 946 5 950
rect 9 946 11 950
rect 15 946 17 950
rect 21 946 23 950
rect 27 946 29 950
rect 33 946 35 950
rect 39 946 41 950
rect 45 946 47 950
rect 51 946 53 950
rect 57 946 59 950
rect 63 946 65 950
rect 69 946 71 950
rect 75 946 77 950
rect 81 946 83 950
rect 87 946 89 950
rect 93 946 95 950
rect 99 946 101 950
rect 105 946 107 950
rect 111 946 113 950
rect 117 946 119 950
rect 123 946 125 950
rect 129 946 131 950
rect 135 946 137 950
rect 141 946 143 950
rect 147 946 149 950
rect 153 946 155 950
rect 159 946 161 950
rect 165 946 167 950
rect 171 946 173 950
rect 177 946 179 950
rect 183 946 185 950
rect 189 946 191 950
rect 195 946 197 950
rect 201 946 203 950
rect 207 946 209 950
rect 213 946 215 950
rect 219 946 221 950
rect 225 946 227 950
rect 231 946 233 950
rect 237 946 239 950
rect 243 946 245 950
rect 249 946 251 950
rect 255 946 257 950
rect 261 946 263 950
rect 267 946 269 950
rect 273 946 275 950
rect 279 946 281 950
rect 285 946 287 950
rect 291 946 293 950
rect 297 946 299 950
rect 303 946 305 950
rect 309 946 311 950
rect 315 946 317 950
rect 321 946 323 950
rect 327 946 329 950
rect 333 946 335 950
rect 339 946 341 950
rect 345 946 347 950
rect 351 946 353 950
rect 357 946 359 950
rect 363 946 365 950
rect 369 946 370 950
rect 2 945 370 946
rect 364 944 370 945
rect 364 940 365 944
rect 369 940 370 944
rect 364 938 370 940
rect 364 934 365 938
rect 369 934 370 938
rect 364 932 370 934
rect 364 928 365 932
rect 369 928 370 932
rect 364 926 370 928
rect 364 922 365 926
rect 369 922 370 926
rect 364 920 370 922
rect 364 916 365 920
rect 369 916 370 920
rect 364 914 370 916
rect 364 910 365 914
rect 369 910 370 914
rect 364 908 370 910
rect 364 904 365 908
rect 369 904 370 908
rect 364 902 370 904
rect 364 898 365 902
rect 369 898 370 902
rect 364 896 370 898
rect 364 892 365 896
rect 369 892 370 896
rect 364 890 370 892
rect 364 886 365 890
rect 369 886 370 890
rect 364 884 370 886
rect 364 880 365 884
rect 369 880 370 884
rect 364 878 370 880
rect 364 874 365 878
rect 369 874 370 878
rect 364 872 370 874
rect 364 868 365 872
rect 369 868 370 872
rect 364 866 370 868
rect 364 862 365 866
rect 369 862 370 866
rect 364 860 370 862
rect 364 856 365 860
rect 369 856 370 860
rect 364 854 370 856
rect 364 850 365 854
rect 369 850 370 854
rect 364 848 370 850
rect 364 844 365 848
rect 369 844 370 848
rect 364 842 370 844
rect 364 838 365 842
rect 369 838 370 842
rect 364 836 370 838
rect 364 832 365 836
rect 369 832 370 836
rect 364 830 370 832
rect 364 826 365 830
rect 369 826 370 830
rect 364 824 370 826
rect 364 820 365 824
rect 369 820 370 824
rect 364 818 370 820
rect 364 814 365 818
rect 369 814 370 818
rect 364 812 370 814
rect 364 808 365 812
rect 369 808 370 812
rect 364 806 370 808
rect 364 802 365 806
rect 369 802 370 806
rect 364 800 370 802
rect 364 796 365 800
rect 369 796 370 800
rect 364 794 370 796
rect 364 790 365 794
rect 369 790 370 794
rect 364 788 370 790
rect 364 784 365 788
rect 369 784 370 788
rect 364 782 370 784
rect 364 778 365 782
rect 369 778 370 782
rect 364 776 370 778
rect 364 772 365 776
rect 369 772 370 776
rect 364 770 370 772
rect 364 766 365 770
rect 369 766 370 770
rect 364 764 370 766
rect 364 760 365 764
rect 369 760 370 764
rect 364 758 370 760
rect 364 754 365 758
rect 369 754 370 758
rect 364 752 370 754
rect 364 748 365 752
rect 369 748 370 752
rect 364 746 370 748
rect 364 742 365 746
rect 369 742 370 746
rect 364 740 370 742
rect 364 736 365 740
rect 369 736 370 740
rect 364 734 370 736
rect 364 730 365 734
rect 369 730 370 734
rect 364 728 370 730
rect 364 724 365 728
rect 369 724 370 728
rect 364 698 370 724
rect 364 694 365 698
rect 369 694 370 698
rect 364 692 370 694
rect 364 688 365 692
rect 369 688 370 692
rect 364 686 370 688
rect 364 682 365 686
rect 369 682 370 686
rect 364 680 370 682
rect 364 676 365 680
rect 369 676 370 680
rect 364 674 370 676
rect 364 670 365 674
rect 369 670 370 674
rect 364 668 370 670
rect 364 664 365 668
rect 369 664 370 668
rect 364 662 370 664
rect 364 658 365 662
rect 369 658 370 662
rect 364 656 370 658
rect 364 652 365 656
rect 369 652 370 656
rect 364 650 370 652
rect 364 646 365 650
rect 369 646 370 650
rect 364 644 370 646
rect 364 640 365 644
rect 369 640 370 644
rect 364 638 370 640
rect 364 634 365 638
rect 369 634 370 638
rect 364 632 370 634
rect 364 628 365 632
rect 369 628 370 632
rect 364 626 370 628
rect 364 622 365 626
rect 369 622 370 626
rect 364 620 370 622
rect 364 616 365 620
rect 369 616 370 620
rect 364 614 370 616
rect 364 610 365 614
rect 369 610 370 614
rect 364 608 370 610
rect 364 604 365 608
rect 369 604 370 608
rect 364 602 370 604
rect 364 598 365 602
rect 369 598 370 602
rect 364 596 370 598
rect 364 592 365 596
rect 369 592 370 596
rect 364 590 370 592
rect 364 586 365 590
rect 369 586 370 590
rect 364 584 370 586
rect 364 580 365 584
rect 369 580 370 584
rect 364 578 370 580
rect 364 574 365 578
rect 369 574 370 578
rect 364 572 370 574
rect 364 568 365 572
rect 369 568 370 572
rect 364 566 370 568
rect 364 562 365 566
rect 369 562 370 566
rect 364 560 370 562
rect 364 556 365 560
rect 369 556 370 560
rect 364 554 370 556
rect 364 550 365 554
rect 369 550 370 554
rect 364 548 370 550
rect 364 544 365 548
rect 369 544 370 548
rect 364 542 370 544
rect 364 538 365 542
rect 369 538 370 542
rect 364 536 370 538
rect 364 532 365 536
rect 369 532 370 536
rect 364 530 370 532
rect 364 526 365 530
rect 369 526 370 530
rect 364 524 370 526
rect 364 520 365 524
rect 369 520 370 524
rect 364 518 370 520
rect 364 514 365 518
rect 369 514 370 518
rect 364 512 370 514
rect 364 508 365 512
rect 369 508 370 512
rect 364 506 370 508
rect 364 502 365 506
rect 369 502 370 506
rect 364 500 370 502
rect 364 496 365 500
rect 369 496 370 500
rect 364 494 370 496
rect 364 490 365 494
rect 369 490 370 494
rect 364 488 370 490
rect 364 484 365 488
rect 369 484 370 488
rect 364 482 370 484
rect 364 478 365 482
rect 369 478 370 482
rect 364 477 370 478
rect 2 476 370 477
rect 2 472 5 476
rect 9 472 11 476
rect 15 472 17 476
rect 21 472 23 476
rect 27 472 29 476
rect 33 472 35 476
rect 39 472 41 476
rect 45 472 47 476
rect 51 472 53 476
rect 57 472 59 476
rect 63 472 65 476
rect 69 472 71 476
rect 75 472 77 476
rect 81 472 83 476
rect 87 472 89 476
rect 93 472 95 476
rect 99 472 101 476
rect 105 472 107 476
rect 111 472 113 476
rect 117 472 119 476
rect 123 472 125 476
rect 129 472 131 476
rect 135 472 137 476
rect 141 472 143 476
rect 147 472 149 476
rect 153 472 155 476
rect 159 472 161 476
rect 165 472 167 476
rect 171 472 173 476
rect 177 472 179 476
rect 183 472 185 476
rect 189 472 191 476
rect 195 472 197 476
rect 201 472 203 476
rect 207 472 209 476
rect 213 472 215 476
rect 219 472 221 476
rect 225 472 227 476
rect 231 472 233 476
rect 237 472 239 476
rect 243 472 245 476
rect 249 472 251 476
rect 255 472 257 476
rect 261 472 263 476
rect 267 472 269 476
rect 273 472 275 476
rect 279 472 281 476
rect 285 472 287 476
rect 291 472 293 476
rect 297 472 299 476
rect 303 472 305 476
rect 309 472 311 476
rect 315 472 317 476
rect 321 472 323 476
rect 327 472 329 476
rect 333 472 335 476
rect 339 472 341 476
rect 345 472 347 476
rect 351 472 353 476
rect 357 472 359 476
rect 363 472 365 476
rect 369 472 370 476
rect 2 471 370 472
rect 364 470 370 471
rect 364 466 365 470
rect 369 466 370 470
rect 364 464 370 466
rect 364 460 365 464
rect 369 460 370 464
rect 364 458 370 460
rect 364 454 365 458
rect 369 454 370 458
rect 364 452 370 454
rect 364 448 365 452
rect 369 448 370 452
rect 364 446 370 448
rect 364 442 365 446
rect 369 442 370 446
rect 364 440 370 442
rect 364 436 365 440
rect 369 436 370 440
rect 364 434 370 436
rect 364 430 365 434
rect 369 430 370 434
rect 364 428 370 430
rect 364 424 365 428
rect 369 424 370 428
rect 364 422 370 424
rect 364 418 365 422
rect 369 418 370 422
rect 364 416 370 418
rect 364 412 365 416
rect 369 412 370 416
rect 364 410 370 412
rect 364 406 365 410
rect 369 406 370 410
rect 364 404 370 406
rect 364 400 365 404
rect 369 400 370 404
rect 364 398 370 400
rect 364 394 365 398
rect 369 394 370 398
rect 364 392 370 394
rect 364 388 365 392
rect 369 388 370 392
rect 364 386 370 388
rect 364 382 365 386
rect 369 382 370 386
rect 364 380 370 382
rect 364 376 365 380
rect 369 376 370 380
rect 364 374 370 376
rect 364 370 365 374
rect 369 370 370 374
rect 364 368 370 370
rect 364 364 365 368
rect 369 364 370 368
rect 364 362 370 364
rect 364 358 365 362
rect 369 358 370 362
rect 364 356 370 358
rect 364 352 365 356
rect 369 352 370 356
rect 364 350 370 352
rect 364 346 365 350
rect 369 346 370 350
rect 364 344 370 346
rect 364 340 365 344
rect 369 340 370 344
rect 364 338 370 340
rect 364 334 365 338
rect 369 334 370 338
rect 364 332 370 334
rect 364 328 365 332
rect 369 328 370 332
rect 364 326 370 328
rect 364 322 365 326
rect 369 322 370 326
rect 364 320 370 322
rect 364 316 365 320
rect 369 316 370 320
rect 364 314 370 316
rect 364 310 365 314
rect 369 310 370 314
rect 364 308 370 310
rect 364 304 365 308
rect 369 304 370 308
rect 364 302 370 304
rect 364 298 365 302
rect 369 298 370 302
rect 364 296 370 298
rect 364 292 365 296
rect 369 292 370 296
rect 364 290 370 292
rect 364 286 365 290
rect 369 286 370 290
rect 364 284 370 286
rect 364 280 365 284
rect 369 280 370 284
rect 364 278 370 280
rect 364 274 365 278
rect 369 274 370 278
rect 364 272 370 274
rect 364 268 365 272
rect 369 268 370 272
rect 364 266 370 268
rect 364 262 365 266
rect 369 262 370 266
rect 364 260 370 262
rect 364 256 365 260
rect 369 256 370 260
rect 364 254 370 256
rect 364 250 365 254
rect 369 250 370 254
rect 364 224 370 250
rect 364 220 365 224
rect 369 220 370 224
rect 364 218 370 220
rect 364 214 365 218
rect 369 214 370 218
rect 364 212 370 214
rect 364 208 365 212
rect 369 208 370 212
rect 364 206 370 208
rect 364 202 365 206
rect 369 202 370 206
rect 364 200 370 202
rect 364 196 365 200
rect 369 196 370 200
rect 364 194 370 196
rect 364 190 365 194
rect 369 190 370 194
rect 364 188 370 190
rect 364 184 365 188
rect 369 184 370 188
rect 364 182 370 184
rect 364 178 365 182
rect 369 178 370 182
rect 364 176 370 178
rect 364 172 365 176
rect 369 172 370 176
rect 364 170 370 172
rect 364 166 365 170
rect 369 166 370 170
rect 364 164 370 166
rect 364 160 365 164
rect 369 160 370 164
rect 364 158 370 160
rect 364 154 365 158
rect 369 154 370 158
rect 364 152 370 154
rect 364 148 365 152
rect 369 148 370 152
rect 364 146 370 148
rect 364 142 365 146
rect 369 142 370 146
rect 364 140 370 142
rect 364 136 365 140
rect 369 136 370 140
rect 364 134 370 136
rect 364 130 365 134
rect 369 130 370 134
rect 364 128 370 130
rect 364 124 365 128
rect 369 124 370 128
rect 364 122 370 124
rect 364 118 365 122
rect 369 118 370 122
rect 364 116 370 118
rect 364 112 365 116
rect 369 112 370 116
rect 364 110 370 112
rect 364 106 365 110
rect 369 106 370 110
rect 364 104 370 106
rect 364 100 365 104
rect 369 100 370 104
rect 364 98 370 100
rect 364 94 365 98
rect 369 94 370 98
rect 364 92 370 94
rect 364 88 365 92
rect 369 88 370 92
rect 364 86 370 88
rect 364 82 365 86
rect 369 82 370 86
rect 364 80 370 82
rect 364 76 365 80
rect 369 76 370 80
rect 364 74 370 76
rect 364 70 365 74
rect 369 70 370 74
rect 364 68 370 70
rect 364 64 365 68
rect 369 64 370 68
rect 364 62 370 64
rect 364 58 365 62
rect 369 58 370 62
rect 364 56 370 58
rect 364 52 365 56
rect 369 52 370 56
rect 364 50 370 52
rect 364 46 365 50
rect 369 46 370 50
rect 364 44 370 46
rect 364 40 365 44
rect 369 40 370 44
rect 364 38 370 40
rect 364 34 365 38
rect 369 34 370 38
rect 364 32 370 34
rect 364 28 365 32
rect 369 28 370 32
rect 364 26 370 28
rect 364 22 365 26
rect 369 22 370 26
rect 364 20 370 22
rect 364 16 365 20
rect 369 16 370 20
rect 364 14 370 16
rect 364 10 365 14
rect 369 10 370 14
rect 364 8 370 10
rect 364 4 365 8
rect 369 4 370 8
rect 364 3 370 4
<< psubstratepcontact >>
rect 365 4258 369 4262
rect 365 4252 369 4256
rect 365 4246 369 4250
rect 365 4240 369 4244
rect 365 4234 369 4238
rect 365 4228 369 4232
rect 365 4222 369 4226
rect 365 4216 369 4220
rect 365 4210 369 4214
rect 365 4204 369 4208
rect 365 4198 369 4202
rect 365 4192 369 4196
rect 365 4186 369 4190
rect 365 4180 369 4184
rect 365 4174 369 4178
rect 365 4168 369 4172
rect 365 4162 369 4166
rect 365 4156 369 4160
rect 365 4150 369 4154
rect 365 4144 369 4148
rect 365 4138 369 4142
rect 365 4132 369 4136
rect 365 4126 369 4130
rect 365 4120 369 4124
rect 365 4114 369 4118
rect 365 4108 369 4112
rect 365 4102 369 4106
rect 365 4096 369 4100
rect 365 4090 369 4094
rect 365 4084 369 4088
rect 365 4078 369 4082
rect 365 4072 369 4076
rect 365 4066 369 4070
rect 365 4060 369 4064
rect 365 4054 369 4058
rect 365 4048 369 4052
rect 365 4042 369 4046
rect 365 4012 369 4016
rect 365 4006 369 4010
rect 365 4000 369 4004
rect 365 3994 369 3998
rect 365 3988 369 3992
rect 365 3982 369 3986
rect 365 3976 369 3980
rect 365 3970 369 3974
rect 365 3964 369 3968
rect 365 3958 369 3962
rect 365 3952 369 3956
rect 365 3946 369 3950
rect 365 3940 369 3944
rect 365 3934 369 3938
rect 365 3928 369 3932
rect 365 3922 369 3926
rect 365 3916 369 3920
rect 365 3910 369 3914
rect 365 3904 369 3908
rect 365 3898 369 3902
rect 365 3892 369 3896
rect 365 3886 369 3890
rect 365 3880 369 3884
rect 365 3874 369 3878
rect 365 3868 369 3872
rect 365 3862 369 3866
rect 365 3856 369 3860
rect 365 3850 369 3854
rect 365 3844 369 3848
rect 365 3838 369 3842
rect 365 3832 369 3836
rect 365 3826 369 3830
rect 365 3820 369 3824
rect 365 3814 369 3818
rect 365 3808 369 3812
rect 365 3802 369 3806
rect 365 3796 369 3800
rect 5 3790 9 3794
rect 11 3790 15 3794
rect 17 3790 21 3794
rect 23 3790 27 3794
rect 29 3790 33 3794
rect 35 3790 39 3794
rect 41 3790 45 3794
rect 47 3790 51 3794
rect 53 3790 57 3794
rect 59 3790 63 3794
rect 65 3790 69 3794
rect 71 3790 75 3794
rect 77 3790 81 3794
rect 83 3790 87 3794
rect 89 3790 93 3794
rect 95 3790 99 3794
rect 101 3790 105 3794
rect 107 3790 111 3794
rect 113 3790 117 3794
rect 119 3790 123 3794
rect 125 3790 129 3794
rect 131 3790 135 3794
rect 137 3790 141 3794
rect 143 3790 147 3794
rect 149 3790 153 3794
rect 155 3790 159 3794
rect 161 3790 165 3794
rect 167 3790 171 3794
rect 173 3790 177 3794
rect 179 3790 183 3794
rect 185 3790 189 3794
rect 191 3790 195 3794
rect 197 3790 201 3794
rect 203 3790 207 3794
rect 209 3790 213 3794
rect 215 3790 219 3794
rect 221 3790 225 3794
rect 227 3790 231 3794
rect 233 3790 237 3794
rect 239 3790 243 3794
rect 245 3790 249 3794
rect 251 3790 255 3794
rect 257 3790 261 3794
rect 263 3790 267 3794
rect 269 3790 273 3794
rect 275 3790 279 3794
rect 281 3790 285 3794
rect 287 3790 291 3794
rect 293 3790 297 3794
rect 299 3790 303 3794
rect 305 3790 309 3794
rect 311 3790 315 3794
rect 317 3790 321 3794
rect 323 3790 327 3794
rect 329 3790 333 3794
rect 335 3790 339 3794
rect 341 3790 345 3794
rect 347 3790 351 3794
rect 353 3790 357 3794
rect 359 3790 363 3794
rect 365 3790 369 3794
rect 365 3784 369 3788
rect 365 3778 369 3782
rect 365 3772 369 3776
rect 365 3766 369 3770
rect 365 3760 369 3764
rect 365 3754 369 3758
rect 365 3748 369 3752
rect 365 3742 369 3746
rect 365 3736 369 3740
rect 365 3730 369 3734
rect 365 3724 369 3728
rect 365 3718 369 3722
rect 365 3712 369 3716
rect 365 3706 369 3710
rect 365 3700 369 3704
rect 365 3694 369 3698
rect 365 3688 369 3692
rect 365 3682 369 3686
rect 365 3676 369 3680
rect 365 3670 369 3674
rect 365 3664 369 3668
rect 365 3658 369 3662
rect 365 3652 369 3656
rect 365 3646 369 3650
rect 365 3640 369 3644
rect 365 3634 369 3638
rect 365 3628 369 3632
rect 365 3622 369 3626
rect 365 3616 369 3620
rect 365 3610 369 3614
rect 365 3604 369 3608
rect 365 3598 369 3602
rect 365 3592 369 3596
rect 365 3586 369 3590
rect 365 3580 369 3584
rect 365 3574 369 3578
rect 365 3568 369 3572
rect 365 3538 369 3542
rect 365 3532 369 3536
rect 365 3526 369 3530
rect 365 3520 369 3524
rect 365 3514 369 3518
rect 365 3508 369 3512
rect 365 3502 369 3506
rect 365 3496 369 3500
rect 365 3490 369 3494
rect 365 3484 369 3488
rect 365 3478 369 3482
rect 365 3472 369 3476
rect 365 3466 369 3470
rect 365 3460 369 3464
rect 365 3454 369 3458
rect 365 3448 369 3452
rect 365 3442 369 3446
rect 365 3436 369 3440
rect 365 3430 369 3434
rect 365 3424 369 3428
rect 365 3418 369 3422
rect 365 3412 369 3416
rect 365 3406 369 3410
rect 365 3400 369 3404
rect 365 3394 369 3398
rect 365 3388 369 3392
rect 365 3382 369 3386
rect 365 3376 369 3380
rect 365 3370 369 3374
rect 365 3364 369 3368
rect 365 3358 369 3362
rect 365 3352 369 3356
rect 365 3346 369 3350
rect 365 3340 369 3344
rect 365 3334 369 3338
rect 365 3328 369 3332
rect 365 3322 369 3326
rect 5 3316 9 3320
rect 11 3316 15 3320
rect 17 3316 21 3320
rect 23 3316 27 3320
rect 29 3316 33 3320
rect 35 3316 39 3320
rect 41 3316 45 3320
rect 47 3316 51 3320
rect 53 3316 57 3320
rect 59 3316 63 3320
rect 65 3316 69 3320
rect 71 3316 75 3320
rect 77 3316 81 3320
rect 83 3316 87 3320
rect 89 3316 93 3320
rect 95 3316 99 3320
rect 101 3316 105 3320
rect 107 3316 111 3320
rect 113 3316 117 3320
rect 119 3316 123 3320
rect 125 3316 129 3320
rect 131 3316 135 3320
rect 137 3316 141 3320
rect 143 3316 147 3320
rect 149 3316 153 3320
rect 155 3316 159 3320
rect 161 3316 165 3320
rect 167 3316 171 3320
rect 173 3316 177 3320
rect 179 3316 183 3320
rect 185 3316 189 3320
rect 191 3316 195 3320
rect 197 3316 201 3320
rect 203 3316 207 3320
rect 209 3316 213 3320
rect 215 3316 219 3320
rect 221 3316 225 3320
rect 227 3316 231 3320
rect 233 3316 237 3320
rect 239 3316 243 3320
rect 245 3316 249 3320
rect 251 3316 255 3320
rect 257 3316 261 3320
rect 263 3316 267 3320
rect 269 3316 273 3320
rect 275 3316 279 3320
rect 281 3316 285 3320
rect 287 3316 291 3320
rect 293 3316 297 3320
rect 299 3316 303 3320
rect 305 3316 309 3320
rect 311 3316 315 3320
rect 317 3316 321 3320
rect 323 3316 327 3320
rect 329 3316 333 3320
rect 335 3316 339 3320
rect 341 3316 345 3320
rect 347 3316 351 3320
rect 353 3316 357 3320
rect 359 3316 363 3320
rect 365 3316 369 3320
rect 365 3310 369 3314
rect 365 3304 369 3308
rect 365 3298 369 3302
rect 365 3292 369 3296
rect 365 3286 369 3290
rect 365 3280 369 3284
rect 365 3274 369 3278
rect 365 3268 369 3272
rect 365 3262 369 3266
rect 365 3256 369 3260
rect 365 3250 369 3254
rect 365 3244 369 3248
rect 365 3238 369 3242
rect 365 3232 369 3236
rect 365 3226 369 3230
rect 365 3220 369 3224
rect 365 3214 369 3218
rect 365 3208 369 3212
rect 365 3202 369 3206
rect 365 3196 369 3200
rect 365 3190 369 3194
rect 365 3184 369 3188
rect 365 3178 369 3182
rect 365 3172 369 3176
rect 365 3166 369 3170
rect 365 3160 369 3164
rect 365 3154 369 3158
rect 365 3148 369 3152
rect 365 3142 369 3146
rect 365 3136 369 3140
rect 365 3130 369 3134
rect 365 3124 369 3128
rect 365 3118 369 3122
rect 365 3112 369 3116
rect 365 3106 369 3110
rect 365 3100 369 3104
rect 365 3094 369 3098
rect 365 3064 369 3068
rect 365 3058 369 3062
rect 365 3052 369 3056
rect 365 3046 369 3050
rect 365 3040 369 3044
rect 365 3034 369 3038
rect 365 3028 369 3032
rect 365 3022 369 3026
rect 365 3016 369 3020
rect 365 3010 369 3014
rect 365 3004 369 3008
rect 365 2998 369 3002
rect 365 2992 369 2996
rect 365 2986 369 2990
rect 365 2980 369 2984
rect 365 2974 369 2978
rect 365 2968 369 2972
rect 365 2962 369 2966
rect 365 2956 369 2960
rect 365 2950 369 2954
rect 365 2944 369 2948
rect 365 2938 369 2942
rect 365 2932 369 2936
rect 365 2926 369 2930
rect 365 2920 369 2924
rect 365 2914 369 2918
rect 365 2908 369 2912
rect 365 2902 369 2906
rect 365 2896 369 2900
rect 365 2890 369 2894
rect 365 2884 369 2888
rect 365 2878 369 2882
rect 365 2872 369 2876
rect 365 2866 369 2870
rect 365 2860 369 2864
rect 365 2854 369 2858
rect 365 2848 369 2852
rect 5 2842 9 2846
rect 11 2842 15 2846
rect 17 2842 21 2846
rect 23 2842 27 2846
rect 29 2842 33 2846
rect 35 2842 39 2846
rect 41 2842 45 2846
rect 47 2842 51 2846
rect 53 2842 57 2846
rect 59 2842 63 2846
rect 65 2842 69 2846
rect 71 2842 75 2846
rect 77 2842 81 2846
rect 83 2842 87 2846
rect 89 2842 93 2846
rect 95 2842 99 2846
rect 101 2842 105 2846
rect 107 2842 111 2846
rect 113 2842 117 2846
rect 119 2842 123 2846
rect 125 2842 129 2846
rect 131 2842 135 2846
rect 137 2842 141 2846
rect 143 2842 147 2846
rect 149 2842 153 2846
rect 155 2842 159 2846
rect 161 2842 165 2846
rect 167 2842 171 2846
rect 173 2842 177 2846
rect 179 2842 183 2846
rect 185 2842 189 2846
rect 191 2842 195 2846
rect 197 2842 201 2846
rect 203 2842 207 2846
rect 209 2842 213 2846
rect 215 2842 219 2846
rect 221 2842 225 2846
rect 227 2842 231 2846
rect 233 2842 237 2846
rect 239 2842 243 2846
rect 245 2842 249 2846
rect 251 2842 255 2846
rect 257 2842 261 2846
rect 263 2842 267 2846
rect 269 2842 273 2846
rect 275 2842 279 2846
rect 281 2842 285 2846
rect 287 2842 291 2846
rect 293 2842 297 2846
rect 299 2842 303 2846
rect 305 2842 309 2846
rect 311 2842 315 2846
rect 317 2842 321 2846
rect 323 2842 327 2846
rect 329 2842 333 2846
rect 335 2842 339 2846
rect 341 2842 345 2846
rect 347 2842 351 2846
rect 353 2842 357 2846
rect 359 2842 363 2846
rect 365 2842 369 2846
rect 365 2836 369 2840
rect 365 2830 369 2834
rect 365 2824 369 2828
rect 365 2818 369 2822
rect 365 2812 369 2816
rect 365 2806 369 2810
rect 365 2800 369 2804
rect 365 2794 369 2798
rect 365 2788 369 2792
rect 365 2782 369 2786
rect 365 2776 369 2780
rect 365 2770 369 2774
rect 365 2764 369 2768
rect 365 2758 369 2762
rect 365 2752 369 2756
rect 365 2746 369 2750
rect 365 2740 369 2744
rect 365 2734 369 2738
rect 365 2728 369 2732
rect 365 2722 369 2726
rect 365 2716 369 2720
rect 365 2710 369 2714
rect 365 2704 369 2708
rect 365 2698 369 2702
rect 365 2692 369 2696
rect 365 2686 369 2690
rect 365 2680 369 2684
rect 365 2674 369 2678
rect 365 2668 369 2672
rect 365 2662 369 2666
rect 365 2656 369 2660
rect 365 2650 369 2654
rect 365 2644 369 2648
rect 365 2638 369 2642
rect 365 2632 369 2636
rect 365 2626 369 2630
rect 365 2620 369 2624
rect 365 2590 369 2594
rect 365 2584 369 2588
rect 365 2578 369 2582
rect 365 2572 369 2576
rect 365 2566 369 2570
rect 365 2560 369 2564
rect 365 2554 369 2558
rect 365 2548 369 2552
rect 365 2542 369 2546
rect 365 2536 369 2540
rect 365 2530 369 2534
rect 365 2524 369 2528
rect 365 2518 369 2522
rect 365 2512 369 2516
rect 365 2506 369 2510
rect 365 2500 369 2504
rect 365 2494 369 2498
rect 365 2488 369 2492
rect 365 2482 369 2486
rect 365 2476 369 2480
rect 365 2470 369 2474
rect 365 2464 369 2468
rect 365 2458 369 2462
rect 365 2452 369 2456
rect 365 2446 369 2450
rect 365 2440 369 2444
rect 365 2434 369 2438
rect 365 2428 369 2432
rect 365 2422 369 2426
rect 365 2416 369 2420
rect 365 2410 369 2414
rect 365 2404 369 2408
rect 365 2398 369 2402
rect 365 2392 369 2396
rect 365 2386 369 2390
rect 365 2380 369 2384
rect 365 2374 369 2378
rect 5 2368 9 2372
rect 11 2368 15 2372
rect 17 2368 21 2372
rect 23 2368 27 2372
rect 29 2368 33 2372
rect 35 2368 39 2372
rect 41 2368 45 2372
rect 47 2368 51 2372
rect 53 2368 57 2372
rect 59 2368 63 2372
rect 65 2368 69 2372
rect 71 2368 75 2372
rect 77 2368 81 2372
rect 83 2368 87 2372
rect 89 2368 93 2372
rect 95 2368 99 2372
rect 101 2368 105 2372
rect 107 2368 111 2372
rect 113 2368 117 2372
rect 119 2368 123 2372
rect 125 2368 129 2372
rect 131 2368 135 2372
rect 137 2368 141 2372
rect 143 2368 147 2372
rect 149 2368 153 2372
rect 155 2368 159 2372
rect 161 2368 165 2372
rect 167 2368 171 2372
rect 173 2368 177 2372
rect 179 2368 183 2372
rect 185 2368 189 2372
rect 191 2368 195 2372
rect 197 2368 201 2372
rect 203 2368 207 2372
rect 209 2368 213 2372
rect 215 2368 219 2372
rect 221 2368 225 2372
rect 227 2368 231 2372
rect 233 2368 237 2372
rect 239 2368 243 2372
rect 245 2368 249 2372
rect 251 2368 255 2372
rect 257 2368 261 2372
rect 263 2368 267 2372
rect 269 2368 273 2372
rect 275 2368 279 2372
rect 281 2368 285 2372
rect 287 2368 291 2372
rect 293 2368 297 2372
rect 299 2368 303 2372
rect 305 2368 309 2372
rect 311 2368 315 2372
rect 317 2368 321 2372
rect 323 2368 327 2372
rect 329 2368 333 2372
rect 335 2368 339 2372
rect 341 2368 345 2372
rect 347 2368 351 2372
rect 353 2368 357 2372
rect 359 2368 363 2372
rect 365 2368 369 2372
rect 365 2362 369 2366
rect 365 2356 369 2360
rect 365 2350 369 2354
rect 365 2344 369 2348
rect 365 2338 369 2342
rect 365 2332 369 2336
rect 365 2326 369 2330
rect 365 2320 369 2324
rect 365 2314 369 2318
rect 365 2308 369 2312
rect 365 2302 369 2306
rect 365 2296 369 2300
rect 365 2290 369 2294
rect 365 2284 369 2288
rect 365 2278 369 2282
rect 365 2272 369 2276
rect 365 2266 369 2270
rect 365 2260 369 2264
rect 365 2254 369 2258
rect 365 2248 369 2252
rect 365 2242 369 2246
rect 365 2236 369 2240
rect 365 2230 369 2234
rect 365 2224 369 2228
rect 365 2218 369 2222
rect 365 2212 369 2216
rect 365 2206 369 2210
rect 365 2200 369 2204
rect 365 2194 369 2198
rect 365 2188 369 2192
rect 365 2182 369 2186
rect 365 2176 369 2180
rect 365 2170 369 2174
rect 365 2164 369 2168
rect 365 2158 369 2162
rect 365 2152 369 2156
rect 365 2146 369 2150
rect 365 2116 369 2120
rect 365 2110 369 2114
rect 365 2104 369 2108
rect 365 2098 369 2102
rect 365 2092 369 2096
rect 365 2086 369 2090
rect 365 2080 369 2084
rect 365 2074 369 2078
rect 365 2068 369 2072
rect 365 2062 369 2066
rect 365 2056 369 2060
rect 365 2050 369 2054
rect 365 2044 369 2048
rect 365 2038 369 2042
rect 365 2032 369 2036
rect 365 2026 369 2030
rect 365 2020 369 2024
rect 365 2014 369 2018
rect 365 2008 369 2012
rect 365 2002 369 2006
rect 365 1996 369 2000
rect 365 1990 369 1994
rect 365 1984 369 1988
rect 365 1978 369 1982
rect 365 1972 369 1976
rect 365 1966 369 1970
rect 365 1960 369 1964
rect 365 1954 369 1958
rect 365 1948 369 1952
rect 365 1942 369 1946
rect 365 1936 369 1940
rect 365 1930 369 1934
rect 365 1924 369 1928
rect 365 1918 369 1922
rect 365 1912 369 1916
rect 365 1906 369 1910
rect 365 1900 369 1904
rect 5 1894 9 1898
rect 11 1894 15 1898
rect 17 1894 21 1898
rect 23 1894 27 1898
rect 29 1894 33 1898
rect 35 1894 39 1898
rect 41 1894 45 1898
rect 47 1894 51 1898
rect 53 1894 57 1898
rect 59 1894 63 1898
rect 65 1894 69 1898
rect 71 1894 75 1898
rect 77 1894 81 1898
rect 83 1894 87 1898
rect 89 1894 93 1898
rect 95 1894 99 1898
rect 101 1894 105 1898
rect 107 1894 111 1898
rect 113 1894 117 1898
rect 119 1894 123 1898
rect 125 1894 129 1898
rect 131 1894 135 1898
rect 137 1894 141 1898
rect 143 1894 147 1898
rect 149 1894 153 1898
rect 155 1894 159 1898
rect 161 1894 165 1898
rect 167 1894 171 1898
rect 173 1894 177 1898
rect 179 1894 183 1898
rect 185 1894 189 1898
rect 191 1894 195 1898
rect 197 1894 201 1898
rect 203 1894 207 1898
rect 209 1894 213 1898
rect 215 1894 219 1898
rect 221 1894 225 1898
rect 227 1894 231 1898
rect 233 1894 237 1898
rect 239 1894 243 1898
rect 245 1894 249 1898
rect 251 1894 255 1898
rect 257 1894 261 1898
rect 263 1894 267 1898
rect 269 1894 273 1898
rect 275 1894 279 1898
rect 281 1894 285 1898
rect 287 1894 291 1898
rect 293 1894 297 1898
rect 299 1894 303 1898
rect 305 1894 309 1898
rect 311 1894 315 1898
rect 317 1894 321 1898
rect 323 1894 327 1898
rect 329 1894 333 1898
rect 335 1894 339 1898
rect 341 1894 345 1898
rect 347 1894 351 1898
rect 353 1894 357 1898
rect 359 1894 363 1898
rect 365 1894 369 1898
rect 365 1888 369 1892
rect 365 1882 369 1886
rect 365 1876 369 1880
rect 365 1870 369 1874
rect 365 1864 369 1868
rect 365 1858 369 1862
rect 365 1852 369 1856
rect 365 1846 369 1850
rect 365 1840 369 1844
rect 365 1834 369 1838
rect 365 1828 369 1832
rect 365 1822 369 1826
rect 365 1816 369 1820
rect 365 1810 369 1814
rect 365 1804 369 1808
rect 365 1798 369 1802
rect 365 1792 369 1796
rect 365 1786 369 1790
rect 365 1780 369 1784
rect 365 1774 369 1778
rect 365 1768 369 1772
rect 365 1762 369 1766
rect 365 1756 369 1760
rect 365 1750 369 1754
rect 365 1744 369 1748
rect 365 1738 369 1742
rect 365 1732 369 1736
rect 365 1726 369 1730
rect 365 1720 369 1724
rect 365 1714 369 1718
rect 365 1708 369 1712
rect 365 1702 369 1706
rect 365 1696 369 1700
rect 365 1690 369 1694
rect 365 1684 369 1688
rect 365 1678 369 1682
rect 365 1672 369 1676
rect 365 1642 369 1646
rect 365 1636 369 1640
rect 365 1630 369 1634
rect 365 1624 369 1628
rect 365 1618 369 1622
rect 365 1612 369 1616
rect 365 1606 369 1610
rect 365 1600 369 1604
rect 365 1594 369 1598
rect 365 1588 369 1592
rect 365 1582 369 1586
rect 365 1576 369 1580
rect 365 1570 369 1574
rect 365 1564 369 1568
rect 365 1558 369 1562
rect 365 1552 369 1556
rect 365 1546 369 1550
rect 365 1540 369 1544
rect 365 1534 369 1538
rect 365 1528 369 1532
rect 365 1522 369 1526
rect 365 1516 369 1520
rect 365 1510 369 1514
rect 365 1504 369 1508
rect 365 1498 369 1502
rect 365 1492 369 1496
rect 365 1486 369 1490
rect 365 1480 369 1484
rect 365 1474 369 1478
rect 365 1468 369 1472
rect 365 1462 369 1466
rect 365 1456 369 1460
rect 365 1450 369 1454
rect 365 1444 369 1448
rect 365 1438 369 1442
rect 365 1432 369 1436
rect 365 1426 369 1430
rect 5 1420 9 1424
rect 11 1420 15 1424
rect 17 1420 21 1424
rect 23 1420 27 1424
rect 29 1420 33 1424
rect 35 1420 39 1424
rect 41 1420 45 1424
rect 47 1420 51 1424
rect 53 1420 57 1424
rect 59 1420 63 1424
rect 65 1420 69 1424
rect 71 1420 75 1424
rect 77 1420 81 1424
rect 83 1420 87 1424
rect 89 1420 93 1424
rect 95 1420 99 1424
rect 101 1420 105 1424
rect 107 1420 111 1424
rect 113 1420 117 1424
rect 119 1420 123 1424
rect 125 1420 129 1424
rect 131 1420 135 1424
rect 137 1420 141 1424
rect 143 1420 147 1424
rect 149 1420 153 1424
rect 155 1420 159 1424
rect 161 1420 165 1424
rect 167 1420 171 1424
rect 173 1420 177 1424
rect 179 1420 183 1424
rect 185 1420 189 1424
rect 191 1420 195 1424
rect 197 1420 201 1424
rect 203 1420 207 1424
rect 209 1420 213 1424
rect 215 1420 219 1424
rect 221 1420 225 1424
rect 227 1420 231 1424
rect 233 1420 237 1424
rect 239 1420 243 1424
rect 245 1420 249 1424
rect 251 1420 255 1424
rect 257 1420 261 1424
rect 263 1420 267 1424
rect 269 1420 273 1424
rect 275 1420 279 1424
rect 281 1420 285 1424
rect 287 1420 291 1424
rect 293 1420 297 1424
rect 299 1420 303 1424
rect 305 1420 309 1424
rect 311 1420 315 1424
rect 317 1420 321 1424
rect 323 1420 327 1424
rect 329 1420 333 1424
rect 335 1420 339 1424
rect 341 1420 345 1424
rect 347 1420 351 1424
rect 353 1420 357 1424
rect 359 1420 363 1424
rect 365 1420 369 1424
rect 365 1414 369 1418
rect 365 1408 369 1412
rect 365 1402 369 1406
rect 365 1396 369 1400
rect 365 1390 369 1394
rect 365 1384 369 1388
rect 365 1378 369 1382
rect 365 1372 369 1376
rect 365 1366 369 1370
rect 365 1360 369 1364
rect 365 1354 369 1358
rect 365 1348 369 1352
rect 365 1342 369 1346
rect 365 1336 369 1340
rect 365 1330 369 1334
rect 365 1324 369 1328
rect 365 1318 369 1322
rect 365 1312 369 1316
rect 365 1306 369 1310
rect 365 1300 369 1304
rect 365 1294 369 1298
rect 365 1288 369 1292
rect 365 1282 369 1286
rect 365 1276 369 1280
rect 365 1270 369 1274
rect 365 1264 369 1268
rect 365 1258 369 1262
rect 365 1252 369 1256
rect 365 1246 369 1250
rect 365 1240 369 1244
rect 365 1234 369 1238
rect 365 1228 369 1232
rect 365 1222 369 1226
rect 365 1216 369 1220
rect 365 1210 369 1214
rect 365 1204 369 1208
rect 365 1198 369 1202
rect 365 1168 369 1172
rect 365 1162 369 1166
rect 365 1156 369 1160
rect 365 1150 369 1154
rect 365 1144 369 1148
rect 365 1138 369 1142
rect 365 1132 369 1136
rect 365 1126 369 1130
rect 365 1120 369 1124
rect 365 1114 369 1118
rect 365 1108 369 1112
rect 365 1102 369 1106
rect 365 1096 369 1100
rect 365 1090 369 1094
rect 365 1084 369 1088
rect 365 1078 369 1082
rect 365 1072 369 1076
rect 365 1066 369 1070
rect 365 1060 369 1064
rect 365 1054 369 1058
rect 365 1048 369 1052
rect 365 1042 369 1046
rect 365 1036 369 1040
rect 365 1030 369 1034
rect 365 1024 369 1028
rect 365 1018 369 1022
rect 365 1012 369 1016
rect 365 1006 369 1010
rect 365 1000 369 1004
rect 365 994 369 998
rect 365 988 369 992
rect 365 982 369 986
rect 365 976 369 980
rect 365 970 369 974
rect 365 964 369 968
rect 365 958 369 962
rect 365 952 369 956
rect 5 946 9 950
rect 11 946 15 950
rect 17 946 21 950
rect 23 946 27 950
rect 29 946 33 950
rect 35 946 39 950
rect 41 946 45 950
rect 47 946 51 950
rect 53 946 57 950
rect 59 946 63 950
rect 65 946 69 950
rect 71 946 75 950
rect 77 946 81 950
rect 83 946 87 950
rect 89 946 93 950
rect 95 946 99 950
rect 101 946 105 950
rect 107 946 111 950
rect 113 946 117 950
rect 119 946 123 950
rect 125 946 129 950
rect 131 946 135 950
rect 137 946 141 950
rect 143 946 147 950
rect 149 946 153 950
rect 155 946 159 950
rect 161 946 165 950
rect 167 946 171 950
rect 173 946 177 950
rect 179 946 183 950
rect 185 946 189 950
rect 191 946 195 950
rect 197 946 201 950
rect 203 946 207 950
rect 209 946 213 950
rect 215 946 219 950
rect 221 946 225 950
rect 227 946 231 950
rect 233 946 237 950
rect 239 946 243 950
rect 245 946 249 950
rect 251 946 255 950
rect 257 946 261 950
rect 263 946 267 950
rect 269 946 273 950
rect 275 946 279 950
rect 281 946 285 950
rect 287 946 291 950
rect 293 946 297 950
rect 299 946 303 950
rect 305 946 309 950
rect 311 946 315 950
rect 317 946 321 950
rect 323 946 327 950
rect 329 946 333 950
rect 335 946 339 950
rect 341 946 345 950
rect 347 946 351 950
rect 353 946 357 950
rect 359 946 363 950
rect 365 946 369 950
rect 365 940 369 944
rect 365 934 369 938
rect 365 928 369 932
rect 365 922 369 926
rect 365 916 369 920
rect 365 910 369 914
rect 365 904 369 908
rect 365 898 369 902
rect 365 892 369 896
rect 365 886 369 890
rect 365 880 369 884
rect 365 874 369 878
rect 365 868 369 872
rect 365 862 369 866
rect 365 856 369 860
rect 365 850 369 854
rect 365 844 369 848
rect 365 838 369 842
rect 365 832 369 836
rect 365 826 369 830
rect 365 820 369 824
rect 365 814 369 818
rect 365 808 369 812
rect 365 802 369 806
rect 365 796 369 800
rect 365 790 369 794
rect 365 784 369 788
rect 365 778 369 782
rect 365 772 369 776
rect 365 766 369 770
rect 365 760 369 764
rect 365 754 369 758
rect 365 748 369 752
rect 365 742 369 746
rect 365 736 369 740
rect 365 730 369 734
rect 365 724 369 728
rect 365 694 369 698
rect 365 688 369 692
rect 365 682 369 686
rect 365 676 369 680
rect 365 670 369 674
rect 365 664 369 668
rect 365 658 369 662
rect 365 652 369 656
rect 365 646 369 650
rect 365 640 369 644
rect 365 634 369 638
rect 365 628 369 632
rect 365 622 369 626
rect 365 616 369 620
rect 365 610 369 614
rect 365 604 369 608
rect 365 598 369 602
rect 365 592 369 596
rect 365 586 369 590
rect 365 580 369 584
rect 365 574 369 578
rect 365 568 369 572
rect 365 562 369 566
rect 365 556 369 560
rect 365 550 369 554
rect 365 544 369 548
rect 365 538 369 542
rect 365 532 369 536
rect 365 526 369 530
rect 365 520 369 524
rect 365 514 369 518
rect 365 508 369 512
rect 365 502 369 506
rect 365 496 369 500
rect 365 490 369 494
rect 365 484 369 488
rect 365 478 369 482
rect 5 472 9 476
rect 11 472 15 476
rect 17 472 21 476
rect 23 472 27 476
rect 29 472 33 476
rect 35 472 39 476
rect 41 472 45 476
rect 47 472 51 476
rect 53 472 57 476
rect 59 472 63 476
rect 65 472 69 476
rect 71 472 75 476
rect 77 472 81 476
rect 83 472 87 476
rect 89 472 93 476
rect 95 472 99 476
rect 101 472 105 476
rect 107 472 111 476
rect 113 472 117 476
rect 119 472 123 476
rect 125 472 129 476
rect 131 472 135 476
rect 137 472 141 476
rect 143 472 147 476
rect 149 472 153 476
rect 155 472 159 476
rect 161 472 165 476
rect 167 472 171 476
rect 173 472 177 476
rect 179 472 183 476
rect 185 472 189 476
rect 191 472 195 476
rect 197 472 201 476
rect 203 472 207 476
rect 209 472 213 476
rect 215 472 219 476
rect 221 472 225 476
rect 227 472 231 476
rect 233 472 237 476
rect 239 472 243 476
rect 245 472 249 476
rect 251 472 255 476
rect 257 472 261 476
rect 263 472 267 476
rect 269 472 273 476
rect 275 472 279 476
rect 281 472 285 476
rect 287 472 291 476
rect 293 472 297 476
rect 299 472 303 476
rect 305 472 309 476
rect 311 472 315 476
rect 317 472 321 476
rect 323 472 327 476
rect 329 472 333 476
rect 335 472 339 476
rect 341 472 345 476
rect 347 472 351 476
rect 353 472 357 476
rect 359 472 363 476
rect 365 472 369 476
rect 365 466 369 470
rect 365 460 369 464
rect 365 454 369 458
rect 365 448 369 452
rect 365 442 369 446
rect 365 436 369 440
rect 365 430 369 434
rect 365 424 369 428
rect 365 418 369 422
rect 365 412 369 416
rect 365 406 369 410
rect 365 400 369 404
rect 365 394 369 398
rect 365 388 369 392
rect 365 382 369 386
rect 365 376 369 380
rect 365 370 369 374
rect 365 364 369 368
rect 365 358 369 362
rect 365 352 369 356
rect 365 346 369 350
rect 365 340 369 344
rect 365 334 369 338
rect 365 328 369 332
rect 365 322 369 326
rect 365 316 369 320
rect 365 310 369 314
rect 365 304 369 308
rect 365 298 369 302
rect 365 292 369 296
rect 365 286 369 290
rect 365 280 369 284
rect 365 274 369 278
rect 365 268 369 272
rect 365 262 369 266
rect 365 256 369 260
rect 365 250 369 254
rect 365 220 369 224
rect 365 214 369 218
rect 365 208 369 212
rect 365 202 369 206
rect 365 196 369 200
rect 365 190 369 194
rect 365 184 369 188
rect 365 178 369 182
rect 365 172 369 176
rect 365 166 369 170
rect 365 160 369 164
rect 365 154 369 158
rect 365 148 369 152
rect 365 142 369 146
rect 365 136 369 140
rect 365 130 369 134
rect 365 124 369 128
rect 365 118 369 122
rect 365 112 369 116
rect 365 106 369 110
rect 365 100 369 104
rect 365 94 369 98
rect 365 88 369 92
rect 365 82 369 86
rect 365 76 369 80
rect 365 70 369 74
rect 365 64 369 68
rect 365 58 369 62
rect 365 52 369 56
rect 365 46 369 50
rect 365 40 369 44
rect 365 34 369 38
rect 365 28 369 32
rect 365 22 369 26
rect 365 16 369 20
rect 365 10 369 14
rect 365 4 369 8
<< polysilicon >>
rect 371 4138 506 4262
rect 371 4134 372 4138
rect 376 4134 506 4138
rect 371 4132 506 4134
rect 371 4128 372 4132
rect 376 4128 506 4132
rect 371 4126 506 4128
rect 371 4122 372 4126
rect 376 4122 506 4126
rect 371 4120 506 4122
rect 371 4116 372 4120
rect 376 4116 506 4120
rect 371 4114 506 4116
rect 371 4110 372 4114
rect 376 4110 506 4114
rect 371 4108 506 4110
rect 371 4104 372 4108
rect 376 4104 506 4108
rect 371 4102 506 4104
rect 371 4098 372 4102
rect 376 4098 506 4102
rect 371 3960 506 4098
rect 371 3956 372 3960
rect 376 3956 501 3960
rect 505 3956 506 3960
rect 371 3954 506 3956
rect 371 3950 372 3954
rect 376 3950 501 3954
rect 505 3950 506 3954
rect 371 3948 506 3950
rect 371 3944 372 3948
rect 376 3944 501 3948
rect 505 3944 506 3948
rect 371 3942 506 3944
rect 371 3938 372 3942
rect 376 3938 501 3942
rect 505 3938 506 3942
rect 371 3936 506 3938
rect 371 3932 372 3936
rect 376 3932 501 3936
rect 505 3932 506 3936
rect 371 3930 506 3932
rect 371 3926 372 3930
rect 376 3926 501 3930
rect 505 3926 506 3930
rect 371 3924 506 3926
rect 371 3920 372 3924
rect 376 3920 501 3924
rect 505 3920 506 3924
rect 371 3664 506 3920
rect 371 3660 372 3664
rect 376 3660 501 3664
rect 505 3660 506 3664
rect 371 3658 506 3660
rect 371 3654 372 3658
rect 376 3654 501 3658
rect 505 3654 506 3658
rect 371 3652 506 3654
rect 371 3648 372 3652
rect 376 3648 501 3652
rect 505 3648 506 3652
rect 371 3646 506 3648
rect 371 3642 372 3646
rect 376 3642 501 3646
rect 505 3642 506 3646
rect 371 3640 506 3642
rect 371 3636 372 3640
rect 376 3636 501 3640
rect 505 3636 506 3640
rect 371 3634 506 3636
rect 371 3630 372 3634
rect 376 3630 501 3634
rect 505 3630 506 3634
rect 371 3628 506 3630
rect 371 3624 372 3628
rect 376 3624 501 3628
rect 505 3624 506 3628
rect 371 3486 506 3624
rect 371 3482 372 3486
rect 376 3482 501 3486
rect 505 3482 506 3486
rect 371 3480 506 3482
rect 371 3476 372 3480
rect 376 3476 501 3480
rect 505 3476 506 3480
rect 371 3474 506 3476
rect 371 3470 372 3474
rect 376 3470 501 3474
rect 505 3470 506 3474
rect 371 3468 506 3470
rect 371 3464 372 3468
rect 376 3464 501 3468
rect 505 3464 506 3468
rect 371 3462 506 3464
rect 371 3458 372 3462
rect 376 3458 501 3462
rect 505 3458 506 3462
rect 371 3456 506 3458
rect 371 3452 372 3456
rect 376 3452 501 3456
rect 505 3452 506 3456
rect 371 3450 506 3452
rect 371 3446 372 3450
rect 376 3446 501 3450
rect 505 3446 506 3450
rect 371 3190 506 3446
rect 371 3186 372 3190
rect 376 3186 501 3190
rect 505 3186 506 3190
rect 371 3184 506 3186
rect 371 3180 372 3184
rect 376 3180 501 3184
rect 505 3180 506 3184
rect 371 3178 506 3180
rect 371 3174 372 3178
rect 376 3174 501 3178
rect 505 3174 506 3178
rect 371 3172 506 3174
rect 371 3168 372 3172
rect 376 3168 501 3172
rect 505 3168 506 3172
rect 371 3166 506 3168
rect 371 3162 372 3166
rect 376 3162 501 3166
rect 505 3162 506 3166
rect 371 3160 506 3162
rect 371 3156 372 3160
rect 376 3156 501 3160
rect 505 3156 506 3160
rect 371 3154 506 3156
rect 371 3150 372 3154
rect 376 3150 501 3154
rect 505 3150 506 3154
rect 371 3012 506 3150
rect 371 3008 372 3012
rect 376 3008 501 3012
rect 505 3008 506 3012
rect 371 3006 506 3008
rect 371 3002 372 3006
rect 376 3002 501 3006
rect 505 3002 506 3006
rect 371 3000 506 3002
rect 371 2996 372 3000
rect 376 2996 501 3000
rect 505 2996 506 3000
rect 371 2994 506 2996
rect 371 2990 372 2994
rect 376 2990 501 2994
rect 505 2990 506 2994
rect 371 2988 506 2990
rect 371 2984 372 2988
rect 376 2984 501 2988
rect 505 2984 506 2988
rect 371 2982 506 2984
rect 371 2978 372 2982
rect 376 2978 501 2982
rect 505 2978 506 2982
rect 371 2976 506 2978
rect 371 2972 372 2976
rect 376 2972 501 2976
rect 505 2972 506 2976
rect 371 2716 506 2972
rect 371 2712 372 2716
rect 376 2712 501 2716
rect 505 2712 506 2716
rect 371 2710 506 2712
rect 371 2706 372 2710
rect 376 2706 501 2710
rect 505 2706 506 2710
rect 371 2704 506 2706
rect 371 2700 372 2704
rect 376 2700 501 2704
rect 505 2700 506 2704
rect 371 2698 506 2700
rect 371 2694 372 2698
rect 376 2694 501 2698
rect 505 2694 506 2698
rect 371 2692 506 2694
rect 371 2688 372 2692
rect 376 2688 501 2692
rect 505 2688 506 2692
rect 371 2686 506 2688
rect 371 2682 372 2686
rect 376 2682 501 2686
rect 505 2682 506 2686
rect 371 2680 506 2682
rect 371 2676 372 2680
rect 376 2676 501 2680
rect 505 2676 506 2680
rect 371 2538 506 2676
rect 371 2534 372 2538
rect 376 2534 501 2538
rect 505 2534 506 2538
rect 371 2532 506 2534
rect 371 2528 372 2532
rect 376 2528 501 2532
rect 505 2528 506 2532
rect 371 2526 506 2528
rect 371 2522 372 2526
rect 376 2522 501 2526
rect 505 2522 506 2526
rect 371 2520 506 2522
rect 371 2516 372 2520
rect 376 2516 501 2520
rect 505 2516 506 2520
rect 371 2514 506 2516
rect 371 2510 372 2514
rect 376 2510 501 2514
rect 505 2510 506 2514
rect 371 2508 506 2510
rect 371 2504 372 2508
rect 376 2504 501 2508
rect 505 2504 506 2508
rect 371 2502 506 2504
rect 371 2498 372 2502
rect 376 2498 501 2502
rect 505 2498 506 2502
rect 371 2242 506 2498
rect 371 2238 372 2242
rect 376 2238 501 2242
rect 505 2238 506 2242
rect 371 2236 506 2238
rect 371 2232 372 2236
rect 376 2232 501 2236
rect 505 2232 506 2236
rect 371 2230 506 2232
rect 371 2226 372 2230
rect 376 2226 501 2230
rect 505 2226 506 2230
rect 371 2224 506 2226
rect 371 2220 372 2224
rect 376 2220 501 2224
rect 505 2220 506 2224
rect 371 2218 506 2220
rect 371 2214 372 2218
rect 376 2214 501 2218
rect 505 2214 506 2218
rect 371 2212 506 2214
rect 371 2208 372 2212
rect 376 2208 501 2212
rect 505 2208 506 2212
rect 371 2206 506 2208
rect 371 2202 372 2206
rect 376 2202 501 2206
rect 505 2202 506 2206
rect 371 2064 506 2202
rect 371 2060 372 2064
rect 376 2060 501 2064
rect 505 2060 506 2064
rect 371 2058 506 2060
rect 371 2054 372 2058
rect 376 2054 501 2058
rect 505 2054 506 2058
rect 371 2052 506 2054
rect 371 2048 372 2052
rect 376 2048 501 2052
rect 505 2048 506 2052
rect 371 2046 506 2048
rect 371 2042 372 2046
rect 376 2042 501 2046
rect 505 2042 506 2046
rect 371 2040 506 2042
rect 371 2036 372 2040
rect 376 2036 501 2040
rect 505 2036 506 2040
rect 371 2034 506 2036
rect 371 2030 372 2034
rect 376 2030 501 2034
rect 505 2030 506 2034
rect 371 2028 506 2030
rect 371 2024 372 2028
rect 376 2024 501 2028
rect 505 2024 506 2028
rect 371 1768 506 2024
rect 371 1764 372 1768
rect 376 1764 501 1768
rect 505 1764 506 1768
rect 371 1762 506 1764
rect 371 1758 372 1762
rect 376 1758 501 1762
rect 505 1758 506 1762
rect 371 1756 506 1758
rect 371 1752 372 1756
rect 376 1752 501 1756
rect 505 1752 506 1756
rect 371 1750 506 1752
rect 371 1746 372 1750
rect 376 1746 501 1750
rect 505 1746 506 1750
rect 371 1744 506 1746
rect 371 1740 372 1744
rect 376 1740 501 1744
rect 505 1740 506 1744
rect 371 1738 506 1740
rect 371 1734 372 1738
rect 376 1734 501 1738
rect 505 1734 506 1738
rect 371 1732 506 1734
rect 371 1728 372 1732
rect 376 1728 501 1732
rect 505 1728 506 1732
rect 371 1590 506 1728
rect 371 1586 372 1590
rect 376 1586 501 1590
rect 505 1586 506 1590
rect 371 1584 506 1586
rect 371 1580 372 1584
rect 376 1580 501 1584
rect 505 1580 506 1584
rect 371 1578 506 1580
rect 371 1574 372 1578
rect 376 1574 501 1578
rect 505 1574 506 1578
rect 371 1572 506 1574
rect 371 1568 372 1572
rect 376 1568 501 1572
rect 505 1568 506 1572
rect 371 1566 506 1568
rect 371 1562 372 1566
rect 376 1562 501 1566
rect 505 1562 506 1566
rect 371 1560 506 1562
rect 371 1556 372 1560
rect 376 1556 501 1560
rect 505 1556 506 1560
rect 371 1554 506 1556
rect 371 1550 372 1554
rect 376 1550 501 1554
rect 505 1550 506 1554
rect 371 1294 506 1550
rect 371 1290 372 1294
rect 376 1290 501 1294
rect 505 1290 506 1294
rect 371 1288 506 1290
rect 371 1284 372 1288
rect 376 1284 501 1288
rect 505 1284 506 1288
rect 371 1282 506 1284
rect 371 1278 372 1282
rect 376 1278 501 1282
rect 505 1278 506 1282
rect 371 1276 506 1278
rect 371 1272 372 1276
rect 376 1272 501 1276
rect 505 1272 506 1276
rect 371 1270 506 1272
rect 371 1266 372 1270
rect 376 1266 501 1270
rect 505 1266 506 1270
rect 371 1264 506 1266
rect 371 1260 372 1264
rect 376 1260 501 1264
rect 505 1260 506 1264
rect 371 1258 506 1260
rect 371 1254 372 1258
rect 376 1254 501 1258
rect 505 1254 506 1258
rect 371 1116 506 1254
rect 371 1112 372 1116
rect 376 1112 501 1116
rect 505 1112 506 1116
rect 371 1110 506 1112
rect 371 1106 372 1110
rect 376 1106 501 1110
rect 505 1106 506 1110
rect 371 1104 506 1106
rect 371 1100 372 1104
rect 376 1100 501 1104
rect 505 1100 506 1104
rect 371 1098 506 1100
rect 371 1094 372 1098
rect 376 1094 501 1098
rect 505 1094 506 1098
rect 371 1092 506 1094
rect 371 1088 372 1092
rect 376 1088 501 1092
rect 505 1088 506 1092
rect 371 1086 506 1088
rect 371 1082 372 1086
rect 376 1082 501 1086
rect 505 1082 506 1086
rect 371 1080 506 1082
rect 371 1076 372 1080
rect 376 1076 501 1080
rect 505 1076 506 1080
rect 371 820 506 1076
rect 371 816 372 820
rect 376 816 501 820
rect 505 816 506 820
rect 371 814 506 816
rect 371 810 372 814
rect 376 810 501 814
rect 505 810 506 814
rect 371 808 506 810
rect 371 804 372 808
rect 376 804 501 808
rect 505 804 506 808
rect 371 802 506 804
rect 371 798 372 802
rect 376 798 501 802
rect 505 798 506 802
rect 371 796 506 798
rect 371 792 372 796
rect 376 792 501 796
rect 505 792 506 796
rect 371 790 506 792
rect 371 786 372 790
rect 376 786 501 790
rect 505 786 506 790
rect 371 784 506 786
rect 371 780 372 784
rect 376 780 501 784
rect 505 780 506 784
rect 371 642 506 780
rect 371 638 372 642
rect 376 638 501 642
rect 505 638 506 642
rect 371 636 506 638
rect 371 632 372 636
rect 376 632 501 636
rect 505 632 506 636
rect 371 630 506 632
rect 371 626 372 630
rect 376 626 501 630
rect 505 626 506 630
rect 371 624 506 626
rect 371 620 372 624
rect 376 620 501 624
rect 505 620 506 624
rect 371 618 506 620
rect 371 614 372 618
rect 376 614 501 618
rect 505 614 506 618
rect 371 612 506 614
rect 371 608 372 612
rect 376 608 501 612
rect 505 608 506 612
rect 371 606 506 608
rect 371 602 372 606
rect 376 602 501 606
rect 505 602 506 606
rect 371 346 506 602
rect 371 342 372 346
rect 376 342 501 346
rect 505 342 506 346
rect 371 340 506 342
rect 371 336 372 340
rect 376 336 501 340
rect 505 336 506 340
rect 371 334 506 336
rect 371 330 372 334
rect 376 330 501 334
rect 505 330 506 334
rect 371 328 506 330
rect 371 324 372 328
rect 376 324 501 328
rect 505 324 506 328
rect 371 322 506 324
rect 371 318 372 322
rect 376 318 501 322
rect 505 318 506 322
rect 371 316 506 318
rect 371 312 372 316
rect 376 312 501 316
rect 505 312 506 316
rect 371 310 506 312
rect 371 306 372 310
rect 376 306 501 310
rect 505 306 506 310
rect 371 168 506 306
rect 371 164 372 168
rect 376 164 506 168
rect 371 162 506 164
rect 371 158 372 162
rect 376 158 506 162
rect 371 156 506 158
rect 371 152 372 156
rect 376 152 506 156
rect 371 150 506 152
rect 371 146 372 150
rect 376 146 506 150
rect 371 144 506 146
rect 371 140 372 144
rect 376 140 506 144
rect 371 138 506 140
rect 371 134 372 138
rect 376 134 506 138
rect 371 132 506 134
rect 371 128 372 132
rect 376 128 506 132
rect 371 4 506 128
<< polycontact >>
rect 372 4134 376 4138
rect 372 4128 376 4132
rect 372 4122 376 4126
rect 372 4116 376 4120
rect 372 4110 376 4114
rect 372 4104 376 4108
rect 372 4098 376 4102
rect 372 3956 376 3960
rect 501 3956 505 3960
rect 372 3950 376 3954
rect 501 3950 505 3954
rect 372 3944 376 3948
rect 501 3944 505 3948
rect 372 3938 376 3942
rect 501 3938 505 3942
rect 372 3932 376 3936
rect 501 3932 505 3936
rect 372 3926 376 3930
rect 501 3926 505 3930
rect 372 3920 376 3924
rect 501 3920 505 3924
rect 372 3660 376 3664
rect 501 3660 505 3664
rect 372 3654 376 3658
rect 501 3654 505 3658
rect 372 3648 376 3652
rect 501 3648 505 3652
rect 372 3642 376 3646
rect 501 3642 505 3646
rect 372 3636 376 3640
rect 501 3636 505 3640
rect 372 3630 376 3634
rect 501 3630 505 3634
rect 372 3624 376 3628
rect 501 3624 505 3628
rect 372 3482 376 3486
rect 501 3482 505 3486
rect 372 3476 376 3480
rect 501 3476 505 3480
rect 372 3470 376 3474
rect 501 3470 505 3474
rect 372 3464 376 3468
rect 501 3464 505 3468
rect 372 3458 376 3462
rect 501 3458 505 3462
rect 372 3452 376 3456
rect 501 3452 505 3456
rect 372 3446 376 3450
rect 501 3446 505 3450
rect 372 3186 376 3190
rect 501 3186 505 3190
rect 372 3180 376 3184
rect 501 3180 505 3184
rect 372 3174 376 3178
rect 501 3174 505 3178
rect 372 3168 376 3172
rect 501 3168 505 3172
rect 372 3162 376 3166
rect 501 3162 505 3166
rect 372 3156 376 3160
rect 501 3156 505 3160
rect 372 3150 376 3154
rect 501 3150 505 3154
rect 372 3008 376 3012
rect 501 3008 505 3012
rect 372 3002 376 3006
rect 501 3002 505 3006
rect 372 2996 376 3000
rect 501 2996 505 3000
rect 372 2990 376 2994
rect 501 2990 505 2994
rect 372 2984 376 2988
rect 501 2984 505 2988
rect 372 2978 376 2982
rect 501 2978 505 2982
rect 372 2972 376 2976
rect 501 2972 505 2976
rect 372 2712 376 2716
rect 501 2712 505 2716
rect 372 2706 376 2710
rect 501 2706 505 2710
rect 372 2700 376 2704
rect 501 2700 505 2704
rect 372 2694 376 2698
rect 501 2694 505 2698
rect 372 2688 376 2692
rect 501 2688 505 2692
rect 372 2682 376 2686
rect 501 2682 505 2686
rect 372 2676 376 2680
rect 501 2676 505 2680
rect 372 2534 376 2538
rect 501 2534 505 2538
rect 372 2528 376 2532
rect 501 2528 505 2532
rect 372 2522 376 2526
rect 501 2522 505 2526
rect 372 2516 376 2520
rect 501 2516 505 2520
rect 372 2510 376 2514
rect 501 2510 505 2514
rect 372 2504 376 2508
rect 501 2504 505 2508
rect 372 2498 376 2502
rect 501 2498 505 2502
rect 372 2238 376 2242
rect 501 2238 505 2242
rect 372 2232 376 2236
rect 501 2232 505 2236
rect 372 2226 376 2230
rect 501 2226 505 2230
rect 372 2220 376 2224
rect 501 2220 505 2224
rect 372 2214 376 2218
rect 501 2214 505 2218
rect 372 2208 376 2212
rect 501 2208 505 2212
rect 372 2202 376 2206
rect 501 2202 505 2206
rect 372 2060 376 2064
rect 501 2060 505 2064
rect 372 2054 376 2058
rect 501 2054 505 2058
rect 372 2048 376 2052
rect 501 2048 505 2052
rect 372 2042 376 2046
rect 501 2042 505 2046
rect 372 2036 376 2040
rect 501 2036 505 2040
rect 372 2030 376 2034
rect 501 2030 505 2034
rect 372 2024 376 2028
rect 501 2024 505 2028
rect 372 1764 376 1768
rect 501 1764 505 1768
rect 372 1758 376 1762
rect 501 1758 505 1762
rect 372 1752 376 1756
rect 501 1752 505 1756
rect 372 1746 376 1750
rect 501 1746 505 1750
rect 372 1740 376 1744
rect 501 1740 505 1744
rect 372 1734 376 1738
rect 501 1734 505 1738
rect 372 1728 376 1732
rect 501 1728 505 1732
rect 372 1586 376 1590
rect 501 1586 505 1590
rect 372 1580 376 1584
rect 501 1580 505 1584
rect 372 1574 376 1578
rect 501 1574 505 1578
rect 372 1568 376 1572
rect 501 1568 505 1572
rect 372 1562 376 1566
rect 501 1562 505 1566
rect 372 1556 376 1560
rect 501 1556 505 1560
rect 372 1550 376 1554
rect 501 1550 505 1554
rect 372 1290 376 1294
rect 501 1290 505 1294
rect 372 1284 376 1288
rect 501 1284 505 1288
rect 372 1278 376 1282
rect 501 1278 505 1282
rect 372 1272 376 1276
rect 501 1272 505 1276
rect 372 1266 376 1270
rect 501 1266 505 1270
rect 372 1260 376 1264
rect 501 1260 505 1264
rect 372 1254 376 1258
rect 501 1254 505 1258
rect 372 1112 376 1116
rect 501 1112 505 1116
rect 372 1106 376 1110
rect 501 1106 505 1110
rect 372 1100 376 1104
rect 501 1100 505 1104
rect 372 1094 376 1098
rect 501 1094 505 1098
rect 372 1088 376 1092
rect 501 1088 505 1092
rect 372 1082 376 1086
rect 501 1082 505 1086
rect 372 1076 376 1080
rect 501 1076 505 1080
rect 372 816 376 820
rect 501 816 505 820
rect 372 810 376 814
rect 501 810 505 814
rect 372 804 376 808
rect 501 804 505 808
rect 372 798 376 802
rect 501 798 505 802
rect 372 792 376 796
rect 501 792 505 796
rect 372 786 376 790
rect 501 786 505 790
rect 372 780 376 784
rect 501 780 505 784
rect 372 638 376 642
rect 501 638 505 642
rect 372 632 376 636
rect 501 632 505 636
rect 372 626 376 630
rect 501 626 505 630
rect 372 620 376 624
rect 501 620 505 624
rect 372 614 376 618
rect 501 614 505 618
rect 372 608 376 612
rect 501 608 505 612
rect 372 602 376 606
rect 501 602 505 606
rect 372 342 376 346
rect 501 342 505 346
rect 372 336 376 340
rect 501 336 505 340
rect 372 330 376 334
rect 501 330 505 334
rect 372 324 376 328
rect 501 324 505 328
rect 372 318 376 322
rect 501 318 505 322
rect 372 312 376 316
rect 501 312 505 316
rect 372 306 376 310
rect 501 306 505 310
rect 372 164 376 168
rect 372 158 376 162
rect 372 152 376 156
rect 372 146 376 150
rect 372 140 376 144
rect 372 134 376 138
rect 372 128 376 132
<< metal1 >>
rect 365 4262 369 4264
rect 365 4256 369 4258
rect 365 4250 369 4252
rect 365 4244 369 4246
rect 365 4238 369 4240
rect 365 4232 369 4234
rect 365 4226 369 4228
rect 365 4220 369 4222
rect 365 4214 369 4216
rect 365 4208 369 4210
rect 365 4202 369 4204
rect 365 4196 369 4198
rect 365 4190 369 4192
rect 365 4184 369 4186
rect 365 4178 369 4180
rect 365 4172 369 4174
rect 365 4166 369 4168
rect 365 4160 369 4162
rect 365 4154 369 4156
rect 365 4148 369 4150
rect 365 4142 369 4144
rect 365 4136 372 4138
rect 369 4134 372 4136
rect 376 4134 412 4138
rect 421 4134 423 4138
rect 427 4134 429 4138
rect 433 4134 435 4138
rect 439 4134 441 4138
rect 450 4134 451 4138
rect 369 4132 451 4134
rect 365 4130 372 4132
rect 369 4128 372 4130
rect 376 4128 412 4132
rect 421 4128 423 4132
rect 427 4128 429 4132
rect 433 4128 435 4132
rect 439 4128 441 4132
rect 450 4128 451 4132
rect 369 4126 451 4128
rect 365 4124 372 4126
rect 369 4122 372 4124
rect 376 4122 412 4126
rect 421 4122 423 4126
rect 427 4122 429 4126
rect 433 4122 435 4126
rect 439 4122 441 4126
rect 450 4122 451 4126
rect 369 4120 451 4122
rect 365 4118 372 4120
rect 369 4116 372 4118
rect 376 4116 412 4120
rect 421 4116 423 4120
rect 427 4116 429 4120
rect 433 4116 435 4120
rect 439 4116 441 4120
rect 450 4116 451 4120
rect 369 4114 451 4116
rect 365 4112 372 4114
rect 369 4110 372 4112
rect 376 4110 412 4114
rect 421 4110 423 4114
rect 427 4110 429 4114
rect 433 4110 435 4114
rect 439 4110 441 4114
rect 450 4110 451 4114
rect 369 4108 451 4110
rect 365 4106 372 4108
rect 369 4104 372 4106
rect 376 4104 412 4108
rect 421 4104 423 4108
rect 427 4104 429 4108
rect 433 4104 435 4108
rect 439 4104 441 4108
rect 450 4104 451 4108
rect 369 4102 451 4104
rect 365 4100 372 4102
rect 369 4098 372 4100
rect 376 4098 412 4102
rect 421 4098 423 4102
rect 427 4098 429 4102
rect 433 4098 435 4102
rect 439 4098 441 4102
rect 450 4098 451 4102
rect 365 4094 369 4096
rect 365 4088 369 4090
rect 388 4090 390 4094
rect 394 4090 397 4094
rect 401 4090 402 4094
rect 384 4088 406 4090
rect 365 4082 369 4084
rect 365 4076 369 4078
rect 365 4070 369 4072
rect 365 4064 369 4066
rect 365 4058 369 4060
rect 382 4084 384 4088
rect 388 4084 390 4088
rect 394 4084 397 4088
rect 401 4084 402 4088
rect 378 4082 406 4084
rect 382 4078 384 4082
rect 388 4078 390 4082
rect 394 4078 397 4082
rect 401 4078 402 4082
rect 378 4076 406 4078
rect 382 4072 384 4076
rect 388 4072 390 4076
rect 394 4072 397 4076
rect 401 4072 402 4076
rect 378 4070 406 4072
rect 382 4066 384 4070
rect 388 4066 390 4070
rect 394 4066 397 4070
rect 401 4066 402 4070
rect 378 4064 406 4066
rect 413 4093 466 4094
rect 413 4089 414 4093
rect 418 4089 420 4093
rect 424 4089 427 4093
rect 431 4089 433 4093
rect 437 4089 439 4093
rect 443 4089 445 4093
rect 449 4090 466 4093
rect 470 4090 471 4094
rect 475 4090 477 4094
rect 481 4090 483 4094
rect 487 4090 489 4094
rect 493 4090 495 4094
rect 499 4090 509 4094
rect 449 4089 513 4090
rect 413 4088 513 4089
rect 413 4087 466 4088
rect 413 4083 414 4087
rect 418 4083 420 4087
rect 424 4083 427 4087
rect 431 4083 433 4087
rect 437 4083 439 4087
rect 443 4083 445 4087
rect 449 4084 466 4087
rect 470 4084 471 4088
rect 475 4084 477 4088
rect 481 4084 483 4088
rect 487 4084 489 4088
rect 493 4084 495 4088
rect 499 4084 509 4088
rect 449 4083 513 4084
rect 413 4082 513 4083
rect 413 4081 466 4082
rect 413 4077 414 4081
rect 418 4077 420 4081
rect 424 4077 427 4081
rect 431 4077 433 4081
rect 437 4077 439 4081
rect 443 4077 445 4081
rect 449 4078 466 4081
rect 470 4078 471 4082
rect 475 4078 477 4082
rect 481 4078 483 4082
rect 487 4078 489 4082
rect 493 4078 495 4082
rect 499 4078 509 4082
rect 449 4077 513 4078
rect 413 4076 513 4077
rect 413 4075 466 4076
rect 413 4071 414 4075
rect 418 4071 420 4075
rect 424 4071 427 4075
rect 431 4071 433 4075
rect 437 4071 439 4075
rect 443 4071 445 4075
rect 449 4072 466 4075
rect 470 4072 471 4076
rect 475 4072 477 4076
rect 481 4072 483 4076
rect 487 4072 489 4076
rect 493 4072 495 4076
rect 499 4072 509 4076
rect 449 4071 513 4072
rect 413 4070 513 4071
rect 413 4069 466 4070
rect 413 4065 414 4069
rect 418 4065 420 4069
rect 424 4065 427 4069
rect 431 4065 433 4069
rect 437 4065 439 4069
rect 443 4065 445 4069
rect 449 4066 466 4069
rect 470 4066 471 4070
rect 475 4066 477 4070
rect 481 4066 483 4070
rect 487 4066 489 4070
rect 493 4066 495 4070
rect 499 4066 509 4070
rect 449 4065 513 4066
rect 413 4064 513 4065
rect 382 4060 384 4064
rect 388 4060 390 4064
rect 394 4060 397 4064
rect 401 4060 402 4064
rect 465 4060 466 4064
rect 470 4060 471 4064
rect 475 4060 477 4064
rect 481 4060 483 4064
rect 487 4060 489 4064
rect 493 4060 495 4064
rect 499 4060 509 4064
rect 378 4058 406 4060
rect 382 4054 384 4058
rect 388 4054 390 4058
rect 394 4054 397 4058
rect 401 4054 402 4058
rect 455 4056 456 4060
rect 460 4056 461 4060
rect 455 4055 461 4056
rect 365 4052 369 4054
rect 365 4046 369 4048
rect 455 4051 456 4055
rect 460 4051 461 4055
rect 465 4058 513 4060
rect 465 4054 466 4058
rect 470 4054 471 4058
rect 475 4054 477 4058
rect 481 4054 483 4058
rect 487 4054 489 4058
rect 493 4054 495 4058
rect 499 4054 509 4058
rect 455 4050 461 4051
rect 455 4046 456 4050
rect 460 4046 509 4050
rect 455 4045 509 4046
rect 455 4041 456 4045
rect 460 4041 509 4045
rect 365 4010 369 4012
rect 365 4004 369 4006
rect 455 4013 456 4017
rect 460 4013 509 4017
rect 455 4012 509 4013
rect 455 4008 456 4012
rect 460 4008 509 4012
rect 455 4007 461 4008
rect 365 3998 369 4000
rect 365 3992 369 3994
rect 365 3986 369 3988
rect 365 3980 369 3982
rect 365 3974 369 3976
rect 382 4000 384 4004
rect 388 4000 390 4004
rect 394 4000 397 4004
rect 401 4000 402 4004
rect 378 3998 406 4000
rect 455 4003 456 4007
rect 460 4003 461 4007
rect 455 4002 461 4003
rect 455 3998 456 4002
rect 460 3998 461 4002
rect 465 4000 466 4004
rect 470 4000 471 4004
rect 475 4000 477 4004
rect 481 4000 483 4004
rect 487 4000 489 4004
rect 493 4000 495 4004
rect 499 4000 509 4004
rect 465 3998 513 4000
rect 382 3994 384 3998
rect 388 3994 390 3998
rect 394 3994 397 3998
rect 401 3994 402 3998
rect 465 3994 466 3998
rect 470 3994 471 3998
rect 475 3994 477 3998
rect 481 3994 483 3998
rect 487 3994 489 3998
rect 493 3994 495 3998
rect 499 3994 509 3998
rect 378 3992 406 3994
rect 382 3988 384 3992
rect 388 3988 390 3992
rect 394 3988 397 3992
rect 401 3988 402 3992
rect 378 3986 406 3988
rect 382 3982 384 3986
rect 388 3982 390 3986
rect 394 3982 397 3986
rect 401 3982 402 3986
rect 378 3980 406 3982
rect 382 3976 384 3980
rect 388 3976 390 3980
rect 394 3976 397 3980
rect 401 3976 402 3980
rect 378 3974 406 3976
rect 382 3970 384 3974
rect 388 3970 390 3974
rect 394 3970 397 3974
rect 401 3970 402 3974
rect 365 3968 369 3970
rect 384 3968 406 3970
rect 388 3964 390 3968
rect 394 3964 397 3968
rect 401 3964 402 3968
rect 413 3993 513 3994
rect 413 3989 414 3993
rect 418 3989 420 3993
rect 424 3989 427 3993
rect 431 3989 433 3993
rect 437 3989 439 3993
rect 443 3989 445 3993
rect 449 3992 513 3993
rect 449 3989 466 3992
rect 413 3988 466 3989
rect 470 3988 471 3992
rect 475 3988 477 3992
rect 481 3988 483 3992
rect 487 3988 489 3992
rect 493 3988 495 3992
rect 499 3988 509 3992
rect 413 3987 513 3988
rect 413 3983 414 3987
rect 418 3983 420 3987
rect 424 3983 427 3987
rect 431 3983 433 3987
rect 437 3983 439 3987
rect 443 3983 445 3987
rect 449 3986 513 3987
rect 449 3983 466 3986
rect 413 3982 466 3983
rect 470 3982 471 3986
rect 475 3982 477 3986
rect 481 3982 483 3986
rect 487 3982 489 3986
rect 493 3982 495 3986
rect 499 3982 509 3986
rect 413 3981 513 3982
rect 413 3977 414 3981
rect 418 3977 420 3981
rect 424 3977 427 3981
rect 431 3977 433 3981
rect 437 3977 439 3981
rect 443 3977 445 3981
rect 449 3980 513 3981
rect 449 3977 466 3980
rect 413 3976 466 3977
rect 470 3976 471 3980
rect 475 3976 477 3980
rect 481 3976 483 3980
rect 487 3976 489 3980
rect 493 3976 495 3980
rect 499 3976 509 3980
rect 413 3975 513 3976
rect 413 3971 414 3975
rect 418 3971 420 3975
rect 424 3971 427 3975
rect 431 3971 433 3975
rect 437 3971 439 3975
rect 443 3971 445 3975
rect 449 3974 513 3975
rect 449 3971 466 3974
rect 413 3970 466 3971
rect 470 3970 471 3974
rect 475 3970 477 3974
rect 481 3970 483 3974
rect 487 3970 489 3974
rect 493 3970 495 3974
rect 499 3970 509 3974
rect 413 3969 513 3970
rect 413 3965 414 3969
rect 418 3965 420 3969
rect 424 3965 427 3969
rect 431 3965 433 3969
rect 437 3965 439 3969
rect 443 3965 445 3969
rect 449 3968 513 3969
rect 449 3965 466 3968
rect 413 3964 466 3965
rect 470 3964 471 3968
rect 475 3964 477 3968
rect 481 3964 483 3968
rect 487 3964 489 3968
rect 493 3964 509 3968
rect 365 3962 369 3964
rect 369 3958 372 3960
rect 365 3956 372 3958
rect 376 3956 412 3960
rect 421 3956 423 3960
rect 427 3956 429 3960
rect 433 3956 435 3960
rect 439 3956 441 3960
rect 450 3956 501 3960
rect 505 3956 509 3960
rect 369 3954 513 3956
rect 369 3952 372 3954
rect 365 3950 372 3952
rect 376 3950 412 3954
rect 421 3950 423 3954
rect 427 3950 429 3954
rect 433 3950 435 3954
rect 439 3950 441 3954
rect 450 3950 501 3954
rect 505 3950 509 3954
rect 369 3948 513 3950
rect 369 3946 372 3948
rect 365 3944 372 3946
rect 376 3944 412 3948
rect 421 3944 423 3948
rect 427 3944 429 3948
rect 433 3944 435 3948
rect 439 3944 441 3948
rect 450 3944 501 3948
rect 505 3944 509 3948
rect 369 3942 513 3944
rect 369 3940 372 3942
rect 365 3938 372 3940
rect 376 3938 412 3942
rect 421 3938 423 3942
rect 427 3938 429 3942
rect 433 3938 435 3942
rect 439 3938 441 3942
rect 450 3938 501 3942
rect 505 3938 509 3942
rect 369 3936 513 3938
rect 369 3934 372 3936
rect 365 3932 372 3934
rect 376 3932 412 3936
rect 421 3932 423 3936
rect 427 3932 429 3936
rect 433 3932 435 3936
rect 439 3932 441 3936
rect 450 3932 501 3936
rect 505 3932 509 3936
rect 369 3930 513 3932
rect 369 3928 372 3930
rect 365 3926 372 3928
rect 376 3926 412 3930
rect 421 3926 423 3930
rect 427 3926 429 3930
rect 433 3926 435 3930
rect 439 3926 441 3930
rect 450 3926 501 3930
rect 505 3926 509 3930
rect 369 3924 513 3926
rect 369 3922 372 3924
rect 365 3920 372 3922
rect 376 3920 412 3924
rect 421 3920 423 3924
rect 427 3920 429 3924
rect 433 3920 435 3924
rect 439 3920 441 3924
rect 450 3920 501 3924
rect 505 3920 509 3924
rect 365 3914 369 3916
rect 365 3908 369 3910
rect 365 3902 369 3904
rect 365 3896 369 3898
rect 365 3890 369 3892
rect 365 3884 369 3886
rect 365 3878 369 3880
rect 365 3872 369 3874
rect 365 3866 369 3868
rect 365 3860 369 3862
rect 365 3854 369 3856
rect 365 3848 369 3850
rect 365 3842 369 3844
rect 365 3836 369 3838
rect 365 3830 369 3832
rect 365 3824 369 3826
rect 365 3818 369 3820
rect 365 3812 369 3814
rect 365 3806 369 3808
rect 365 3800 369 3802
rect 365 3794 369 3796
rect 3 3790 5 3794
rect 9 3790 11 3794
rect 15 3790 17 3794
rect 21 3790 23 3794
rect 27 3790 29 3794
rect 33 3790 35 3794
rect 39 3790 41 3794
rect 45 3790 47 3794
rect 51 3790 53 3794
rect 57 3790 59 3794
rect 63 3790 65 3794
rect 69 3790 71 3794
rect 75 3790 77 3794
rect 81 3790 83 3794
rect 87 3790 89 3794
rect 93 3790 95 3794
rect 99 3790 101 3794
rect 105 3790 107 3794
rect 111 3790 113 3794
rect 117 3790 119 3794
rect 123 3790 125 3794
rect 129 3790 131 3794
rect 135 3790 137 3794
rect 141 3790 143 3794
rect 147 3790 149 3794
rect 153 3790 155 3794
rect 159 3790 161 3794
rect 165 3790 167 3794
rect 171 3790 173 3794
rect 177 3790 179 3794
rect 183 3790 185 3794
rect 189 3790 191 3794
rect 195 3790 197 3794
rect 201 3790 203 3794
rect 207 3790 209 3794
rect 213 3790 215 3794
rect 219 3790 221 3794
rect 225 3790 227 3794
rect 231 3790 233 3794
rect 237 3790 239 3794
rect 243 3790 245 3794
rect 249 3790 251 3794
rect 255 3790 257 3794
rect 261 3790 263 3794
rect 267 3790 269 3794
rect 273 3790 275 3794
rect 279 3790 281 3794
rect 285 3790 287 3794
rect 291 3790 293 3794
rect 297 3790 299 3794
rect 303 3790 305 3794
rect 309 3790 311 3794
rect 315 3790 317 3794
rect 321 3790 323 3794
rect 327 3790 329 3794
rect 333 3790 335 3794
rect 339 3790 341 3794
rect 345 3790 347 3794
rect 351 3790 353 3794
rect 357 3790 359 3794
rect 363 3790 365 3794
rect 365 3788 369 3790
rect 365 3782 369 3784
rect 365 3776 369 3778
rect 365 3770 369 3772
rect 365 3764 369 3766
rect 365 3758 369 3760
rect 365 3752 369 3754
rect 365 3746 369 3748
rect 365 3740 369 3742
rect 365 3734 369 3736
rect 365 3728 369 3730
rect 365 3722 369 3724
rect 365 3716 369 3718
rect 365 3710 369 3712
rect 365 3704 369 3706
rect 365 3698 369 3700
rect 365 3692 369 3694
rect 365 3686 369 3688
rect 365 3680 369 3682
rect 365 3674 369 3676
rect 365 3668 369 3670
rect 365 3662 372 3664
rect 369 3660 372 3662
rect 376 3660 412 3664
rect 421 3660 423 3664
rect 427 3660 429 3664
rect 433 3660 435 3664
rect 439 3660 441 3664
rect 450 3660 501 3664
rect 505 3660 509 3664
rect 369 3658 513 3660
rect 365 3656 372 3658
rect 369 3654 372 3656
rect 376 3654 412 3658
rect 421 3654 423 3658
rect 427 3654 429 3658
rect 433 3654 435 3658
rect 439 3654 441 3658
rect 450 3654 501 3658
rect 505 3654 509 3658
rect 369 3652 513 3654
rect 365 3650 372 3652
rect 369 3648 372 3650
rect 376 3648 412 3652
rect 421 3648 423 3652
rect 427 3648 429 3652
rect 433 3648 435 3652
rect 439 3648 441 3652
rect 450 3648 501 3652
rect 505 3648 509 3652
rect 369 3646 513 3648
rect 365 3644 372 3646
rect 369 3642 372 3644
rect 376 3642 412 3646
rect 421 3642 423 3646
rect 427 3642 429 3646
rect 433 3642 435 3646
rect 439 3642 441 3646
rect 450 3642 501 3646
rect 505 3642 509 3646
rect 369 3640 513 3642
rect 365 3638 372 3640
rect 369 3636 372 3638
rect 376 3636 412 3640
rect 421 3636 423 3640
rect 427 3636 429 3640
rect 433 3636 435 3640
rect 439 3636 441 3640
rect 450 3636 501 3640
rect 505 3636 509 3640
rect 369 3634 513 3636
rect 365 3632 372 3634
rect 369 3630 372 3632
rect 376 3630 412 3634
rect 421 3630 423 3634
rect 427 3630 429 3634
rect 433 3630 435 3634
rect 439 3630 441 3634
rect 450 3630 501 3634
rect 505 3630 509 3634
rect 369 3628 513 3630
rect 365 3626 372 3628
rect 369 3624 372 3626
rect 376 3624 412 3628
rect 421 3624 423 3628
rect 427 3624 429 3628
rect 433 3624 435 3628
rect 439 3624 441 3628
rect 450 3624 501 3628
rect 505 3624 509 3628
rect 365 3620 369 3622
rect 365 3614 369 3616
rect 388 3616 390 3620
rect 394 3616 397 3620
rect 401 3616 402 3620
rect 384 3614 406 3616
rect 365 3608 369 3610
rect 365 3602 369 3604
rect 365 3596 369 3598
rect 365 3590 369 3592
rect 365 3584 369 3586
rect 382 3610 384 3614
rect 388 3610 390 3614
rect 394 3610 397 3614
rect 401 3610 402 3614
rect 378 3608 406 3610
rect 382 3604 384 3608
rect 388 3604 390 3608
rect 394 3604 397 3608
rect 401 3604 402 3608
rect 378 3602 406 3604
rect 382 3598 384 3602
rect 388 3598 390 3602
rect 394 3598 397 3602
rect 401 3598 402 3602
rect 378 3596 406 3598
rect 382 3592 384 3596
rect 388 3592 390 3596
rect 394 3592 397 3596
rect 401 3592 402 3596
rect 378 3590 406 3592
rect 413 3619 465 3620
rect 413 3615 414 3619
rect 418 3615 420 3619
rect 424 3615 427 3619
rect 431 3615 433 3619
rect 437 3615 439 3619
rect 443 3615 445 3619
rect 449 3616 465 3619
rect 469 3616 471 3620
rect 475 3616 477 3620
rect 481 3616 483 3620
rect 487 3616 489 3620
rect 493 3616 509 3620
rect 449 3615 513 3616
rect 413 3614 513 3615
rect 413 3613 465 3614
rect 413 3609 414 3613
rect 418 3609 420 3613
rect 424 3609 427 3613
rect 431 3609 433 3613
rect 437 3609 439 3613
rect 443 3609 445 3613
rect 449 3610 465 3613
rect 469 3610 471 3614
rect 475 3610 477 3614
rect 481 3610 483 3614
rect 487 3610 489 3614
rect 493 3610 495 3614
rect 499 3610 509 3614
rect 449 3609 513 3610
rect 413 3608 513 3609
rect 413 3607 465 3608
rect 413 3603 414 3607
rect 418 3603 420 3607
rect 424 3603 427 3607
rect 431 3603 433 3607
rect 437 3603 439 3607
rect 443 3603 445 3607
rect 449 3604 465 3607
rect 469 3604 471 3608
rect 475 3604 477 3608
rect 481 3604 483 3608
rect 487 3604 489 3608
rect 493 3604 495 3608
rect 499 3604 509 3608
rect 449 3603 513 3604
rect 413 3602 513 3603
rect 413 3601 465 3602
rect 413 3597 414 3601
rect 418 3597 420 3601
rect 424 3597 427 3601
rect 431 3597 433 3601
rect 437 3597 439 3601
rect 443 3597 445 3601
rect 449 3598 465 3601
rect 469 3598 471 3602
rect 475 3598 477 3602
rect 481 3598 483 3602
rect 487 3598 489 3602
rect 493 3598 495 3602
rect 499 3598 509 3602
rect 449 3597 513 3598
rect 413 3596 513 3597
rect 413 3595 465 3596
rect 413 3591 414 3595
rect 418 3591 420 3595
rect 424 3591 427 3595
rect 431 3591 433 3595
rect 437 3591 439 3595
rect 443 3591 445 3595
rect 449 3592 465 3595
rect 469 3592 471 3596
rect 475 3592 477 3596
rect 481 3592 483 3596
rect 487 3592 489 3596
rect 493 3592 495 3596
rect 499 3592 509 3596
rect 449 3591 513 3592
rect 413 3590 513 3591
rect 382 3586 384 3590
rect 388 3586 390 3590
rect 394 3586 397 3590
rect 401 3586 402 3590
rect 469 3586 471 3590
rect 475 3586 477 3590
rect 481 3586 483 3590
rect 487 3586 489 3590
rect 493 3586 495 3590
rect 499 3586 509 3590
rect 378 3584 406 3586
rect 382 3580 384 3584
rect 388 3580 390 3584
rect 394 3580 397 3584
rect 401 3580 402 3584
rect 455 3582 456 3586
rect 460 3582 461 3586
rect 455 3581 461 3582
rect 365 3578 369 3580
rect 365 3572 369 3574
rect 455 3577 456 3581
rect 460 3577 461 3581
rect 465 3584 513 3586
rect 469 3580 471 3584
rect 475 3580 477 3584
rect 481 3580 483 3584
rect 487 3580 489 3584
rect 493 3580 495 3584
rect 499 3580 509 3584
rect 455 3576 461 3577
rect 455 3572 456 3576
rect 460 3572 509 3576
rect 455 3571 509 3572
rect 455 3567 456 3571
rect 460 3567 509 3571
rect 365 3536 369 3538
rect 365 3530 369 3532
rect 455 3539 456 3543
rect 460 3539 509 3543
rect 455 3538 509 3539
rect 455 3534 456 3538
rect 460 3534 509 3538
rect 455 3533 461 3534
rect 365 3524 369 3526
rect 365 3518 369 3520
rect 365 3512 369 3514
rect 365 3506 369 3508
rect 365 3500 369 3502
rect 382 3526 384 3530
rect 388 3526 390 3530
rect 394 3526 397 3530
rect 401 3526 402 3530
rect 378 3524 406 3526
rect 455 3529 456 3533
rect 460 3529 461 3533
rect 455 3528 461 3529
rect 455 3524 456 3528
rect 460 3524 461 3528
rect 469 3526 471 3530
rect 475 3526 477 3530
rect 481 3526 483 3530
rect 487 3526 489 3530
rect 493 3526 495 3530
rect 499 3526 509 3530
rect 465 3524 513 3526
rect 382 3520 384 3524
rect 388 3520 390 3524
rect 394 3520 397 3524
rect 401 3520 402 3524
rect 469 3520 471 3524
rect 475 3520 477 3524
rect 481 3520 483 3524
rect 487 3520 489 3524
rect 493 3520 495 3524
rect 499 3520 509 3524
rect 378 3518 406 3520
rect 382 3514 384 3518
rect 388 3514 390 3518
rect 394 3514 397 3518
rect 401 3514 402 3518
rect 378 3512 406 3514
rect 382 3508 384 3512
rect 388 3508 390 3512
rect 394 3508 397 3512
rect 401 3508 402 3512
rect 378 3506 406 3508
rect 382 3502 384 3506
rect 388 3502 390 3506
rect 394 3502 397 3506
rect 401 3502 402 3506
rect 378 3500 406 3502
rect 382 3496 384 3500
rect 388 3496 390 3500
rect 394 3496 397 3500
rect 401 3496 402 3500
rect 365 3494 369 3496
rect 384 3494 406 3496
rect 388 3490 390 3494
rect 394 3490 397 3494
rect 401 3490 402 3494
rect 413 3519 513 3520
rect 413 3515 414 3519
rect 418 3515 420 3519
rect 424 3515 427 3519
rect 431 3515 433 3519
rect 437 3515 439 3519
rect 443 3515 445 3519
rect 449 3518 513 3519
rect 449 3515 465 3518
rect 413 3514 465 3515
rect 469 3514 471 3518
rect 475 3514 477 3518
rect 481 3514 483 3518
rect 487 3514 489 3518
rect 493 3514 495 3518
rect 499 3514 509 3518
rect 413 3513 513 3514
rect 413 3509 414 3513
rect 418 3509 420 3513
rect 424 3509 427 3513
rect 431 3509 433 3513
rect 437 3509 439 3513
rect 443 3509 445 3513
rect 449 3512 513 3513
rect 449 3509 465 3512
rect 413 3508 465 3509
rect 469 3508 471 3512
rect 475 3508 477 3512
rect 481 3508 483 3512
rect 487 3508 489 3512
rect 493 3508 495 3512
rect 499 3508 509 3512
rect 413 3507 513 3508
rect 413 3503 414 3507
rect 418 3503 420 3507
rect 424 3503 427 3507
rect 431 3503 433 3507
rect 437 3503 439 3507
rect 443 3503 445 3507
rect 449 3506 513 3507
rect 449 3503 465 3506
rect 413 3502 465 3503
rect 469 3502 471 3506
rect 475 3502 477 3506
rect 481 3502 483 3506
rect 487 3502 489 3506
rect 493 3502 495 3506
rect 499 3502 509 3506
rect 413 3501 513 3502
rect 413 3497 414 3501
rect 418 3497 420 3501
rect 424 3497 427 3501
rect 431 3497 433 3501
rect 437 3497 439 3501
rect 443 3497 445 3501
rect 449 3500 513 3501
rect 449 3497 465 3500
rect 413 3496 465 3497
rect 469 3496 471 3500
rect 475 3496 477 3500
rect 481 3496 483 3500
rect 487 3496 489 3500
rect 493 3496 495 3500
rect 499 3496 509 3500
rect 413 3495 513 3496
rect 413 3491 414 3495
rect 418 3491 420 3495
rect 424 3491 427 3495
rect 431 3491 433 3495
rect 437 3491 439 3495
rect 443 3491 445 3495
rect 449 3494 513 3495
rect 449 3491 465 3494
rect 413 3490 465 3491
rect 469 3490 471 3494
rect 475 3490 477 3494
rect 481 3490 483 3494
rect 487 3490 489 3494
rect 493 3490 509 3494
rect 365 3488 369 3490
rect 369 3484 372 3486
rect 365 3482 372 3484
rect 376 3482 412 3486
rect 421 3482 423 3486
rect 427 3482 429 3486
rect 433 3482 435 3486
rect 439 3482 441 3486
rect 450 3482 501 3486
rect 505 3482 509 3486
rect 369 3480 513 3482
rect 369 3478 372 3480
rect 365 3476 372 3478
rect 376 3476 412 3480
rect 421 3476 423 3480
rect 427 3476 429 3480
rect 433 3476 435 3480
rect 439 3476 441 3480
rect 450 3476 501 3480
rect 505 3476 509 3480
rect 369 3474 513 3476
rect 369 3472 372 3474
rect 365 3470 372 3472
rect 376 3470 412 3474
rect 421 3470 423 3474
rect 427 3470 429 3474
rect 433 3470 435 3474
rect 439 3470 441 3474
rect 450 3470 501 3474
rect 505 3470 509 3474
rect 369 3468 513 3470
rect 369 3466 372 3468
rect 365 3464 372 3466
rect 376 3464 412 3468
rect 421 3464 423 3468
rect 427 3464 429 3468
rect 433 3464 435 3468
rect 439 3464 441 3468
rect 450 3464 501 3468
rect 505 3464 509 3468
rect 369 3462 513 3464
rect 369 3460 372 3462
rect 365 3458 372 3460
rect 376 3458 412 3462
rect 421 3458 423 3462
rect 427 3458 429 3462
rect 433 3458 435 3462
rect 439 3458 441 3462
rect 450 3458 501 3462
rect 505 3458 509 3462
rect 369 3456 513 3458
rect 369 3454 372 3456
rect 365 3452 372 3454
rect 376 3452 412 3456
rect 421 3452 423 3456
rect 427 3452 429 3456
rect 433 3452 435 3456
rect 439 3452 441 3456
rect 450 3452 501 3456
rect 505 3452 509 3456
rect 369 3450 513 3452
rect 369 3448 372 3450
rect 365 3446 372 3448
rect 376 3446 412 3450
rect 421 3446 423 3450
rect 427 3446 429 3450
rect 433 3446 435 3450
rect 439 3446 441 3450
rect 450 3446 501 3450
rect 505 3446 509 3450
rect 365 3440 369 3442
rect 365 3434 369 3436
rect 365 3428 369 3430
rect 365 3422 369 3424
rect 365 3416 369 3418
rect 365 3410 369 3412
rect 365 3404 369 3406
rect 365 3398 369 3400
rect 365 3392 369 3394
rect 365 3386 369 3388
rect 365 3380 369 3382
rect 365 3374 369 3376
rect 365 3368 369 3370
rect 365 3362 369 3364
rect 365 3356 369 3358
rect 365 3350 369 3352
rect 365 3344 369 3346
rect 365 3338 369 3340
rect 365 3332 369 3334
rect 365 3326 369 3328
rect 365 3320 369 3322
rect 3 3316 5 3320
rect 9 3316 11 3320
rect 15 3316 17 3320
rect 21 3316 23 3320
rect 27 3316 29 3320
rect 33 3316 35 3320
rect 39 3316 41 3320
rect 45 3316 47 3320
rect 51 3316 53 3320
rect 57 3316 59 3320
rect 63 3316 65 3320
rect 69 3316 71 3320
rect 75 3316 77 3320
rect 81 3316 83 3320
rect 87 3316 89 3320
rect 93 3316 95 3320
rect 99 3316 101 3320
rect 105 3316 107 3320
rect 111 3316 113 3320
rect 117 3316 119 3320
rect 123 3316 125 3320
rect 129 3316 131 3320
rect 135 3316 137 3320
rect 141 3316 143 3320
rect 147 3316 149 3320
rect 153 3316 155 3320
rect 159 3316 161 3320
rect 165 3316 167 3320
rect 171 3316 173 3320
rect 177 3316 179 3320
rect 183 3316 185 3320
rect 189 3316 191 3320
rect 195 3316 197 3320
rect 201 3316 203 3320
rect 207 3316 209 3320
rect 213 3316 215 3320
rect 219 3316 221 3320
rect 225 3316 227 3320
rect 231 3316 233 3320
rect 237 3316 239 3320
rect 243 3316 245 3320
rect 249 3316 251 3320
rect 255 3316 257 3320
rect 261 3316 263 3320
rect 267 3316 269 3320
rect 273 3316 275 3320
rect 279 3316 281 3320
rect 285 3316 287 3320
rect 291 3316 293 3320
rect 297 3316 299 3320
rect 303 3316 305 3320
rect 309 3316 311 3320
rect 315 3316 317 3320
rect 321 3316 323 3320
rect 327 3316 329 3320
rect 333 3316 335 3320
rect 339 3316 341 3320
rect 345 3316 347 3320
rect 351 3316 353 3320
rect 357 3316 359 3320
rect 363 3316 365 3320
rect 365 3314 369 3316
rect 365 3308 369 3310
rect 365 3302 369 3304
rect 365 3296 369 3298
rect 365 3290 369 3292
rect 365 3284 369 3286
rect 365 3278 369 3280
rect 365 3272 369 3274
rect 365 3266 369 3268
rect 365 3260 369 3262
rect 365 3254 369 3256
rect 365 3248 369 3250
rect 365 3242 369 3244
rect 365 3236 369 3238
rect 365 3230 369 3232
rect 365 3224 369 3226
rect 365 3218 369 3220
rect 365 3212 369 3214
rect 365 3206 369 3208
rect 365 3200 369 3202
rect 365 3194 369 3196
rect 365 3188 372 3190
rect 369 3186 372 3188
rect 376 3186 412 3190
rect 421 3186 423 3190
rect 427 3186 429 3190
rect 433 3186 435 3190
rect 439 3186 441 3190
rect 450 3186 501 3190
rect 505 3186 509 3190
rect 369 3184 513 3186
rect 365 3182 372 3184
rect 369 3180 372 3182
rect 376 3180 412 3184
rect 421 3180 423 3184
rect 427 3180 429 3184
rect 433 3180 435 3184
rect 439 3180 441 3184
rect 450 3180 501 3184
rect 505 3180 509 3184
rect 369 3178 513 3180
rect 365 3176 372 3178
rect 369 3174 372 3176
rect 376 3174 412 3178
rect 421 3174 423 3178
rect 427 3174 429 3178
rect 433 3174 435 3178
rect 439 3174 441 3178
rect 450 3174 501 3178
rect 505 3174 509 3178
rect 369 3172 513 3174
rect 365 3170 372 3172
rect 369 3168 372 3170
rect 376 3168 412 3172
rect 421 3168 423 3172
rect 427 3168 429 3172
rect 433 3168 435 3172
rect 439 3168 441 3172
rect 450 3168 501 3172
rect 505 3168 509 3172
rect 369 3166 513 3168
rect 365 3164 372 3166
rect 369 3162 372 3164
rect 376 3162 412 3166
rect 421 3162 423 3166
rect 427 3162 429 3166
rect 433 3162 435 3166
rect 439 3162 441 3166
rect 450 3162 501 3166
rect 505 3162 509 3166
rect 369 3160 513 3162
rect 365 3158 372 3160
rect 369 3156 372 3158
rect 376 3156 412 3160
rect 421 3156 423 3160
rect 427 3156 429 3160
rect 433 3156 435 3160
rect 439 3156 441 3160
rect 450 3156 501 3160
rect 505 3156 509 3160
rect 369 3154 513 3156
rect 365 3152 372 3154
rect 369 3150 372 3152
rect 376 3150 412 3154
rect 421 3150 423 3154
rect 427 3150 429 3154
rect 433 3150 435 3154
rect 439 3150 441 3154
rect 450 3150 501 3154
rect 505 3150 509 3154
rect 365 3146 369 3148
rect 365 3140 369 3142
rect 388 3142 390 3146
rect 394 3142 397 3146
rect 401 3142 402 3146
rect 384 3140 406 3142
rect 365 3134 369 3136
rect 365 3128 369 3130
rect 365 3122 369 3124
rect 365 3116 369 3118
rect 365 3110 369 3112
rect 382 3136 384 3140
rect 388 3136 390 3140
rect 394 3136 397 3140
rect 401 3136 402 3140
rect 378 3134 406 3136
rect 382 3130 384 3134
rect 388 3130 390 3134
rect 394 3130 397 3134
rect 401 3130 402 3134
rect 378 3128 406 3130
rect 382 3124 384 3128
rect 388 3124 390 3128
rect 394 3124 397 3128
rect 401 3124 402 3128
rect 378 3122 406 3124
rect 382 3118 384 3122
rect 388 3118 390 3122
rect 394 3118 397 3122
rect 401 3118 402 3122
rect 378 3116 406 3118
rect 413 3145 465 3146
rect 413 3141 414 3145
rect 418 3141 420 3145
rect 424 3141 427 3145
rect 431 3141 433 3145
rect 437 3141 439 3145
rect 443 3141 445 3145
rect 449 3142 465 3145
rect 469 3142 471 3146
rect 475 3142 477 3146
rect 481 3142 483 3146
rect 487 3142 489 3146
rect 493 3142 509 3146
rect 449 3141 513 3142
rect 413 3140 513 3141
rect 413 3139 465 3140
rect 413 3135 414 3139
rect 418 3135 420 3139
rect 424 3135 427 3139
rect 431 3135 433 3139
rect 437 3135 439 3139
rect 443 3135 445 3139
rect 449 3136 465 3139
rect 469 3136 471 3140
rect 475 3136 477 3140
rect 481 3136 483 3140
rect 487 3136 489 3140
rect 493 3136 495 3140
rect 499 3136 509 3140
rect 449 3135 513 3136
rect 413 3134 513 3135
rect 413 3133 465 3134
rect 413 3129 414 3133
rect 418 3129 420 3133
rect 424 3129 427 3133
rect 431 3129 433 3133
rect 437 3129 439 3133
rect 443 3129 445 3133
rect 449 3130 465 3133
rect 469 3130 471 3134
rect 475 3130 477 3134
rect 481 3130 483 3134
rect 487 3130 489 3134
rect 493 3130 495 3134
rect 499 3130 509 3134
rect 449 3129 513 3130
rect 413 3128 513 3129
rect 413 3127 465 3128
rect 413 3123 414 3127
rect 418 3123 420 3127
rect 424 3123 427 3127
rect 431 3123 433 3127
rect 437 3123 439 3127
rect 443 3123 445 3127
rect 449 3124 465 3127
rect 469 3124 471 3128
rect 475 3124 477 3128
rect 481 3124 483 3128
rect 487 3124 489 3128
rect 493 3124 495 3128
rect 499 3124 509 3128
rect 449 3123 513 3124
rect 413 3122 513 3123
rect 413 3121 465 3122
rect 413 3117 414 3121
rect 418 3117 420 3121
rect 424 3117 427 3121
rect 431 3117 433 3121
rect 437 3117 439 3121
rect 443 3117 445 3121
rect 449 3118 465 3121
rect 469 3118 471 3122
rect 475 3118 477 3122
rect 481 3118 483 3122
rect 487 3118 489 3122
rect 493 3118 495 3122
rect 499 3118 509 3122
rect 449 3117 513 3118
rect 413 3116 513 3117
rect 382 3112 384 3116
rect 388 3112 390 3116
rect 394 3112 397 3116
rect 401 3112 402 3116
rect 469 3112 471 3116
rect 475 3112 477 3116
rect 481 3112 483 3116
rect 487 3112 489 3116
rect 493 3112 495 3116
rect 499 3112 509 3116
rect 378 3110 406 3112
rect 382 3106 384 3110
rect 388 3106 390 3110
rect 394 3106 397 3110
rect 401 3106 402 3110
rect 455 3108 456 3112
rect 460 3108 461 3112
rect 455 3107 461 3108
rect 365 3104 369 3106
rect 365 3098 369 3100
rect 455 3103 456 3107
rect 460 3103 461 3107
rect 465 3110 513 3112
rect 469 3106 471 3110
rect 475 3106 477 3110
rect 481 3106 483 3110
rect 487 3106 489 3110
rect 493 3106 495 3110
rect 499 3106 509 3110
rect 455 3102 461 3103
rect 455 3098 456 3102
rect 460 3098 509 3102
rect 455 3097 509 3098
rect 455 3093 456 3097
rect 460 3093 509 3097
rect 365 3062 369 3064
rect 365 3056 369 3058
rect 455 3065 456 3069
rect 460 3065 509 3069
rect 455 3064 509 3065
rect 455 3060 456 3064
rect 460 3060 509 3064
rect 455 3059 461 3060
rect 365 3050 369 3052
rect 365 3044 369 3046
rect 365 3038 369 3040
rect 365 3032 369 3034
rect 365 3026 369 3028
rect 382 3052 384 3056
rect 388 3052 390 3056
rect 394 3052 397 3056
rect 401 3052 402 3056
rect 378 3050 406 3052
rect 455 3055 456 3059
rect 460 3055 461 3059
rect 455 3054 461 3055
rect 455 3050 456 3054
rect 460 3050 461 3054
rect 469 3052 471 3056
rect 475 3052 477 3056
rect 481 3052 483 3056
rect 487 3052 489 3056
rect 493 3052 495 3056
rect 499 3052 509 3056
rect 465 3050 513 3052
rect 382 3046 384 3050
rect 388 3046 390 3050
rect 394 3046 397 3050
rect 401 3046 402 3050
rect 469 3046 471 3050
rect 475 3046 477 3050
rect 481 3046 483 3050
rect 487 3046 489 3050
rect 493 3046 495 3050
rect 499 3046 509 3050
rect 378 3044 406 3046
rect 382 3040 384 3044
rect 388 3040 390 3044
rect 394 3040 397 3044
rect 401 3040 402 3044
rect 378 3038 406 3040
rect 382 3034 384 3038
rect 388 3034 390 3038
rect 394 3034 397 3038
rect 401 3034 402 3038
rect 378 3032 406 3034
rect 382 3028 384 3032
rect 388 3028 390 3032
rect 394 3028 397 3032
rect 401 3028 402 3032
rect 378 3026 406 3028
rect 382 3022 384 3026
rect 388 3022 390 3026
rect 394 3022 397 3026
rect 401 3022 402 3026
rect 365 3020 369 3022
rect 384 3020 406 3022
rect 388 3016 390 3020
rect 394 3016 397 3020
rect 401 3016 402 3020
rect 413 3045 513 3046
rect 413 3041 414 3045
rect 418 3041 420 3045
rect 424 3041 427 3045
rect 431 3041 433 3045
rect 437 3041 439 3045
rect 443 3041 445 3045
rect 449 3044 513 3045
rect 449 3041 465 3044
rect 413 3040 465 3041
rect 469 3040 471 3044
rect 475 3040 477 3044
rect 481 3040 483 3044
rect 487 3040 489 3044
rect 493 3040 495 3044
rect 499 3040 509 3044
rect 413 3039 513 3040
rect 413 3035 414 3039
rect 418 3035 420 3039
rect 424 3035 427 3039
rect 431 3035 433 3039
rect 437 3035 439 3039
rect 443 3035 445 3039
rect 449 3038 513 3039
rect 449 3035 465 3038
rect 413 3034 465 3035
rect 469 3034 471 3038
rect 475 3034 477 3038
rect 481 3034 483 3038
rect 487 3034 489 3038
rect 493 3034 495 3038
rect 499 3034 509 3038
rect 413 3033 513 3034
rect 413 3029 414 3033
rect 418 3029 420 3033
rect 424 3029 427 3033
rect 431 3029 433 3033
rect 437 3029 439 3033
rect 443 3029 445 3033
rect 449 3032 513 3033
rect 449 3029 465 3032
rect 413 3028 465 3029
rect 469 3028 471 3032
rect 475 3028 477 3032
rect 481 3028 483 3032
rect 487 3028 489 3032
rect 493 3028 495 3032
rect 499 3028 509 3032
rect 413 3027 513 3028
rect 413 3023 414 3027
rect 418 3023 420 3027
rect 424 3023 427 3027
rect 431 3023 433 3027
rect 437 3023 439 3027
rect 443 3023 445 3027
rect 449 3026 513 3027
rect 449 3023 465 3026
rect 413 3022 465 3023
rect 469 3022 471 3026
rect 475 3022 477 3026
rect 481 3022 483 3026
rect 487 3022 489 3026
rect 493 3022 495 3026
rect 499 3022 509 3026
rect 413 3021 513 3022
rect 413 3017 414 3021
rect 418 3017 420 3021
rect 424 3017 427 3021
rect 431 3017 433 3021
rect 437 3017 439 3021
rect 443 3017 445 3021
rect 449 3020 513 3021
rect 449 3017 465 3020
rect 413 3016 465 3017
rect 469 3016 471 3020
rect 475 3016 477 3020
rect 481 3016 483 3020
rect 487 3016 489 3020
rect 493 3016 509 3020
rect 365 3014 369 3016
rect 369 3010 372 3012
rect 365 3008 372 3010
rect 376 3008 412 3012
rect 421 3008 423 3012
rect 427 3008 429 3012
rect 433 3008 435 3012
rect 439 3008 441 3012
rect 450 3008 501 3012
rect 505 3008 509 3012
rect 369 3006 513 3008
rect 369 3004 372 3006
rect 365 3002 372 3004
rect 376 3002 412 3006
rect 421 3002 423 3006
rect 427 3002 429 3006
rect 433 3002 435 3006
rect 439 3002 441 3006
rect 450 3002 501 3006
rect 505 3002 509 3006
rect 369 3000 513 3002
rect 369 2998 372 3000
rect 365 2996 372 2998
rect 376 2996 412 3000
rect 421 2996 423 3000
rect 427 2996 429 3000
rect 433 2996 435 3000
rect 439 2996 441 3000
rect 450 2996 501 3000
rect 505 2996 509 3000
rect 369 2994 513 2996
rect 369 2992 372 2994
rect 365 2990 372 2992
rect 376 2990 412 2994
rect 421 2990 423 2994
rect 427 2990 429 2994
rect 433 2990 435 2994
rect 439 2990 441 2994
rect 450 2990 501 2994
rect 505 2990 509 2994
rect 369 2988 513 2990
rect 369 2986 372 2988
rect 365 2984 372 2986
rect 376 2984 412 2988
rect 421 2984 423 2988
rect 427 2984 429 2988
rect 433 2984 435 2988
rect 439 2984 441 2988
rect 450 2984 501 2988
rect 505 2984 509 2988
rect 369 2982 513 2984
rect 369 2980 372 2982
rect 365 2978 372 2980
rect 376 2978 412 2982
rect 421 2978 423 2982
rect 427 2978 429 2982
rect 433 2978 435 2982
rect 439 2978 441 2982
rect 450 2978 501 2982
rect 505 2978 509 2982
rect 369 2976 513 2978
rect 369 2974 372 2976
rect 365 2972 372 2974
rect 376 2972 412 2976
rect 421 2972 423 2976
rect 427 2972 429 2976
rect 433 2972 435 2976
rect 439 2972 441 2976
rect 450 2972 501 2976
rect 505 2972 509 2976
rect 365 2966 369 2968
rect 365 2960 369 2962
rect 365 2954 369 2956
rect 365 2948 369 2950
rect 365 2942 369 2944
rect 365 2936 369 2938
rect 365 2930 369 2932
rect 365 2924 369 2926
rect 365 2918 369 2920
rect 365 2912 369 2914
rect 365 2906 369 2908
rect 365 2900 369 2902
rect 365 2894 369 2896
rect 365 2888 369 2890
rect 365 2882 369 2884
rect 365 2876 369 2878
rect 365 2870 369 2872
rect 365 2864 369 2866
rect 365 2858 369 2860
rect 365 2852 369 2854
rect 365 2846 369 2848
rect 3 2842 5 2846
rect 9 2842 11 2846
rect 15 2842 17 2846
rect 21 2842 23 2846
rect 27 2842 29 2846
rect 33 2842 35 2846
rect 39 2842 41 2846
rect 45 2842 47 2846
rect 51 2842 53 2846
rect 57 2842 59 2846
rect 63 2842 65 2846
rect 69 2842 71 2846
rect 75 2842 77 2846
rect 81 2842 83 2846
rect 87 2842 89 2846
rect 93 2842 95 2846
rect 99 2842 101 2846
rect 105 2842 107 2846
rect 111 2842 113 2846
rect 117 2842 119 2846
rect 123 2842 125 2846
rect 129 2842 131 2846
rect 135 2842 137 2846
rect 141 2842 143 2846
rect 147 2842 149 2846
rect 153 2842 155 2846
rect 159 2842 161 2846
rect 165 2842 167 2846
rect 171 2842 173 2846
rect 177 2842 179 2846
rect 183 2842 185 2846
rect 189 2842 191 2846
rect 195 2842 197 2846
rect 201 2842 203 2846
rect 207 2842 209 2846
rect 213 2842 215 2846
rect 219 2842 221 2846
rect 225 2842 227 2846
rect 231 2842 233 2846
rect 237 2842 239 2846
rect 243 2842 245 2846
rect 249 2842 251 2846
rect 255 2842 257 2846
rect 261 2842 263 2846
rect 267 2842 269 2846
rect 273 2842 275 2846
rect 279 2842 281 2846
rect 285 2842 287 2846
rect 291 2842 293 2846
rect 297 2842 299 2846
rect 303 2842 305 2846
rect 309 2842 311 2846
rect 315 2842 317 2846
rect 321 2842 323 2846
rect 327 2842 329 2846
rect 333 2842 335 2846
rect 339 2842 341 2846
rect 345 2842 347 2846
rect 351 2842 353 2846
rect 357 2842 359 2846
rect 363 2842 365 2846
rect 365 2840 369 2842
rect 365 2834 369 2836
rect 365 2828 369 2830
rect 365 2822 369 2824
rect 365 2816 369 2818
rect 365 2810 369 2812
rect 365 2804 369 2806
rect 365 2798 369 2800
rect 365 2792 369 2794
rect 365 2786 369 2788
rect 365 2780 369 2782
rect 365 2774 369 2776
rect 365 2768 369 2770
rect 365 2762 369 2764
rect 365 2756 369 2758
rect 365 2750 369 2752
rect 365 2744 369 2746
rect 365 2738 369 2740
rect 365 2732 369 2734
rect 365 2726 369 2728
rect 365 2720 369 2722
rect 365 2714 372 2716
rect 369 2712 372 2714
rect 376 2712 412 2716
rect 421 2712 423 2716
rect 427 2712 429 2716
rect 433 2712 435 2716
rect 439 2712 441 2716
rect 450 2712 501 2716
rect 505 2712 509 2716
rect 369 2710 513 2712
rect 365 2708 372 2710
rect 369 2706 372 2708
rect 376 2706 412 2710
rect 421 2706 423 2710
rect 427 2706 429 2710
rect 433 2706 435 2710
rect 439 2706 441 2710
rect 450 2706 501 2710
rect 505 2706 509 2710
rect 369 2704 513 2706
rect 365 2702 372 2704
rect 369 2700 372 2702
rect 376 2700 412 2704
rect 421 2700 423 2704
rect 427 2700 429 2704
rect 433 2700 435 2704
rect 439 2700 441 2704
rect 450 2700 501 2704
rect 505 2700 509 2704
rect 369 2698 513 2700
rect 365 2696 372 2698
rect 369 2694 372 2696
rect 376 2694 412 2698
rect 421 2694 423 2698
rect 427 2694 429 2698
rect 433 2694 435 2698
rect 439 2694 441 2698
rect 450 2694 501 2698
rect 505 2694 509 2698
rect 369 2692 513 2694
rect 365 2690 372 2692
rect 369 2688 372 2690
rect 376 2688 412 2692
rect 421 2688 423 2692
rect 427 2688 429 2692
rect 433 2688 435 2692
rect 439 2688 441 2692
rect 450 2688 501 2692
rect 505 2688 509 2692
rect 369 2686 513 2688
rect 365 2684 372 2686
rect 369 2682 372 2684
rect 376 2682 412 2686
rect 421 2682 423 2686
rect 427 2682 429 2686
rect 433 2682 435 2686
rect 439 2682 441 2686
rect 450 2682 501 2686
rect 505 2682 509 2686
rect 369 2680 513 2682
rect 365 2678 372 2680
rect 369 2676 372 2678
rect 376 2676 412 2680
rect 421 2676 423 2680
rect 427 2676 429 2680
rect 433 2676 435 2680
rect 439 2676 441 2680
rect 450 2676 501 2680
rect 505 2676 509 2680
rect 365 2672 369 2674
rect 365 2666 369 2668
rect 388 2668 390 2672
rect 394 2668 397 2672
rect 401 2668 402 2672
rect 384 2666 406 2668
rect 365 2660 369 2662
rect 365 2654 369 2656
rect 365 2648 369 2650
rect 365 2642 369 2644
rect 365 2636 369 2638
rect 382 2662 384 2666
rect 388 2662 390 2666
rect 394 2662 397 2666
rect 401 2662 402 2666
rect 378 2660 406 2662
rect 382 2656 384 2660
rect 388 2656 390 2660
rect 394 2656 397 2660
rect 401 2656 402 2660
rect 378 2654 406 2656
rect 382 2650 384 2654
rect 388 2650 390 2654
rect 394 2650 397 2654
rect 401 2650 402 2654
rect 378 2648 406 2650
rect 382 2644 384 2648
rect 388 2644 390 2648
rect 394 2644 397 2648
rect 401 2644 402 2648
rect 378 2642 406 2644
rect 413 2671 465 2672
rect 413 2667 414 2671
rect 418 2667 420 2671
rect 424 2667 427 2671
rect 431 2667 433 2671
rect 437 2667 439 2671
rect 443 2667 445 2671
rect 449 2668 465 2671
rect 469 2668 471 2672
rect 475 2668 477 2672
rect 481 2668 483 2672
rect 487 2668 489 2672
rect 493 2668 509 2672
rect 449 2667 513 2668
rect 413 2666 513 2667
rect 413 2665 465 2666
rect 413 2661 414 2665
rect 418 2661 420 2665
rect 424 2661 427 2665
rect 431 2661 433 2665
rect 437 2661 439 2665
rect 443 2661 445 2665
rect 449 2662 465 2665
rect 469 2662 471 2666
rect 475 2662 477 2666
rect 481 2662 483 2666
rect 487 2662 489 2666
rect 493 2662 495 2666
rect 499 2662 509 2666
rect 449 2661 513 2662
rect 413 2660 513 2661
rect 413 2659 465 2660
rect 413 2655 414 2659
rect 418 2655 420 2659
rect 424 2655 427 2659
rect 431 2655 433 2659
rect 437 2655 439 2659
rect 443 2655 445 2659
rect 449 2656 465 2659
rect 469 2656 471 2660
rect 475 2656 477 2660
rect 481 2656 483 2660
rect 487 2656 489 2660
rect 493 2656 495 2660
rect 499 2656 509 2660
rect 449 2655 513 2656
rect 413 2654 513 2655
rect 413 2653 465 2654
rect 413 2649 414 2653
rect 418 2649 420 2653
rect 424 2649 427 2653
rect 431 2649 433 2653
rect 437 2649 439 2653
rect 443 2649 445 2653
rect 449 2650 465 2653
rect 469 2650 471 2654
rect 475 2650 477 2654
rect 481 2650 483 2654
rect 487 2650 489 2654
rect 493 2650 495 2654
rect 499 2650 509 2654
rect 449 2649 513 2650
rect 413 2648 513 2649
rect 413 2647 465 2648
rect 413 2643 414 2647
rect 418 2643 420 2647
rect 424 2643 427 2647
rect 431 2643 433 2647
rect 437 2643 439 2647
rect 443 2643 445 2647
rect 449 2644 465 2647
rect 469 2644 471 2648
rect 475 2644 477 2648
rect 481 2644 483 2648
rect 487 2644 489 2648
rect 493 2644 495 2648
rect 499 2644 509 2648
rect 449 2643 513 2644
rect 413 2642 513 2643
rect 382 2638 384 2642
rect 388 2638 390 2642
rect 394 2638 397 2642
rect 401 2638 402 2642
rect 469 2638 471 2642
rect 475 2638 477 2642
rect 481 2638 483 2642
rect 487 2638 489 2642
rect 493 2638 495 2642
rect 499 2638 509 2642
rect 378 2636 406 2638
rect 382 2632 384 2636
rect 388 2632 390 2636
rect 394 2632 397 2636
rect 401 2632 402 2636
rect 455 2634 456 2638
rect 460 2634 461 2638
rect 455 2633 461 2634
rect 365 2630 369 2632
rect 365 2624 369 2626
rect 455 2629 456 2633
rect 460 2629 461 2633
rect 465 2636 513 2638
rect 469 2632 471 2636
rect 475 2632 477 2636
rect 481 2632 483 2636
rect 487 2632 489 2636
rect 493 2632 495 2636
rect 499 2632 509 2636
rect 455 2628 461 2629
rect 455 2624 456 2628
rect 460 2624 509 2628
rect 455 2623 509 2624
rect 455 2619 456 2623
rect 460 2619 509 2623
rect 365 2588 369 2590
rect 365 2582 369 2584
rect 455 2591 456 2595
rect 460 2591 509 2595
rect 455 2590 509 2591
rect 455 2586 456 2590
rect 460 2586 509 2590
rect 455 2585 461 2586
rect 365 2576 369 2578
rect 365 2570 369 2572
rect 365 2564 369 2566
rect 365 2558 369 2560
rect 365 2552 369 2554
rect 382 2578 384 2582
rect 388 2578 390 2582
rect 394 2578 397 2582
rect 401 2578 402 2582
rect 378 2576 406 2578
rect 455 2581 456 2585
rect 460 2581 461 2585
rect 455 2580 461 2581
rect 455 2576 456 2580
rect 460 2576 461 2580
rect 469 2578 471 2582
rect 475 2578 477 2582
rect 481 2578 483 2582
rect 487 2578 489 2582
rect 493 2578 495 2582
rect 499 2578 509 2582
rect 465 2576 513 2578
rect 382 2572 384 2576
rect 388 2572 390 2576
rect 394 2572 397 2576
rect 401 2572 402 2576
rect 469 2572 471 2576
rect 475 2572 477 2576
rect 481 2572 483 2576
rect 487 2572 489 2576
rect 493 2572 495 2576
rect 499 2572 509 2576
rect 378 2570 406 2572
rect 382 2566 384 2570
rect 388 2566 390 2570
rect 394 2566 397 2570
rect 401 2566 402 2570
rect 378 2564 406 2566
rect 382 2560 384 2564
rect 388 2560 390 2564
rect 394 2560 397 2564
rect 401 2560 402 2564
rect 378 2558 406 2560
rect 382 2554 384 2558
rect 388 2554 390 2558
rect 394 2554 397 2558
rect 401 2554 402 2558
rect 378 2552 406 2554
rect 382 2548 384 2552
rect 388 2548 390 2552
rect 394 2548 397 2552
rect 401 2548 402 2552
rect 365 2546 369 2548
rect 384 2546 406 2548
rect 388 2542 390 2546
rect 394 2542 397 2546
rect 401 2542 402 2546
rect 413 2571 513 2572
rect 413 2567 414 2571
rect 418 2567 420 2571
rect 424 2567 427 2571
rect 431 2567 433 2571
rect 437 2567 439 2571
rect 443 2567 445 2571
rect 449 2570 513 2571
rect 449 2567 465 2570
rect 413 2566 465 2567
rect 469 2566 471 2570
rect 475 2566 477 2570
rect 481 2566 483 2570
rect 487 2566 489 2570
rect 493 2566 495 2570
rect 499 2566 509 2570
rect 413 2565 513 2566
rect 413 2561 414 2565
rect 418 2561 420 2565
rect 424 2561 427 2565
rect 431 2561 433 2565
rect 437 2561 439 2565
rect 443 2561 445 2565
rect 449 2564 513 2565
rect 449 2561 465 2564
rect 413 2560 465 2561
rect 469 2560 471 2564
rect 475 2560 477 2564
rect 481 2560 483 2564
rect 487 2560 489 2564
rect 493 2560 495 2564
rect 499 2560 509 2564
rect 413 2559 513 2560
rect 413 2555 414 2559
rect 418 2555 420 2559
rect 424 2555 427 2559
rect 431 2555 433 2559
rect 437 2555 439 2559
rect 443 2555 445 2559
rect 449 2558 513 2559
rect 449 2555 465 2558
rect 413 2554 465 2555
rect 469 2554 471 2558
rect 475 2554 477 2558
rect 481 2554 483 2558
rect 487 2554 489 2558
rect 493 2554 495 2558
rect 499 2554 509 2558
rect 413 2553 513 2554
rect 413 2549 414 2553
rect 418 2549 420 2553
rect 424 2549 427 2553
rect 431 2549 433 2553
rect 437 2549 439 2553
rect 443 2549 445 2553
rect 449 2552 513 2553
rect 449 2549 465 2552
rect 413 2548 465 2549
rect 469 2548 471 2552
rect 475 2548 477 2552
rect 481 2548 483 2552
rect 487 2548 489 2552
rect 493 2548 495 2552
rect 499 2548 509 2552
rect 413 2547 513 2548
rect 413 2543 414 2547
rect 418 2543 420 2547
rect 424 2543 427 2547
rect 431 2543 433 2547
rect 437 2543 439 2547
rect 443 2543 445 2547
rect 449 2546 513 2547
rect 449 2543 465 2546
rect 413 2542 465 2543
rect 469 2542 471 2546
rect 475 2542 477 2546
rect 481 2542 483 2546
rect 487 2542 489 2546
rect 493 2542 509 2546
rect 365 2540 369 2542
rect 369 2536 372 2538
rect 365 2534 372 2536
rect 376 2534 412 2538
rect 421 2534 423 2538
rect 427 2534 429 2538
rect 433 2534 435 2538
rect 439 2534 441 2538
rect 450 2534 501 2538
rect 505 2534 509 2538
rect 369 2532 513 2534
rect 369 2530 372 2532
rect 365 2528 372 2530
rect 376 2528 412 2532
rect 421 2528 423 2532
rect 427 2528 429 2532
rect 433 2528 435 2532
rect 439 2528 441 2532
rect 450 2528 501 2532
rect 505 2528 509 2532
rect 369 2526 513 2528
rect 369 2524 372 2526
rect 365 2522 372 2524
rect 376 2522 412 2526
rect 421 2522 423 2526
rect 427 2522 429 2526
rect 433 2522 435 2526
rect 439 2522 441 2526
rect 450 2522 501 2526
rect 505 2522 509 2526
rect 369 2520 513 2522
rect 369 2518 372 2520
rect 365 2516 372 2518
rect 376 2516 412 2520
rect 421 2516 423 2520
rect 427 2516 429 2520
rect 433 2516 435 2520
rect 439 2516 441 2520
rect 450 2516 501 2520
rect 505 2516 509 2520
rect 369 2514 513 2516
rect 369 2512 372 2514
rect 365 2510 372 2512
rect 376 2510 412 2514
rect 421 2510 423 2514
rect 427 2510 429 2514
rect 433 2510 435 2514
rect 439 2510 441 2514
rect 450 2510 501 2514
rect 505 2510 509 2514
rect 369 2508 513 2510
rect 369 2506 372 2508
rect 365 2504 372 2506
rect 376 2504 412 2508
rect 421 2504 423 2508
rect 427 2504 429 2508
rect 433 2504 435 2508
rect 439 2504 441 2508
rect 450 2504 501 2508
rect 505 2504 509 2508
rect 369 2502 513 2504
rect 369 2500 372 2502
rect 365 2498 372 2500
rect 376 2498 412 2502
rect 421 2498 423 2502
rect 427 2498 429 2502
rect 433 2498 435 2502
rect 439 2498 441 2502
rect 450 2498 501 2502
rect 505 2498 509 2502
rect 365 2492 369 2494
rect 365 2486 369 2488
rect 365 2480 369 2482
rect 365 2474 369 2476
rect 365 2468 369 2470
rect 365 2462 369 2464
rect 365 2456 369 2458
rect 365 2450 369 2452
rect 365 2444 369 2446
rect 365 2438 369 2440
rect 365 2432 369 2434
rect 365 2426 369 2428
rect 365 2420 369 2422
rect 365 2414 369 2416
rect 365 2408 369 2410
rect 365 2402 369 2404
rect 365 2396 369 2398
rect 365 2390 369 2392
rect 365 2384 369 2386
rect 365 2378 369 2380
rect 365 2372 369 2374
rect 3 2368 5 2372
rect 9 2368 11 2372
rect 15 2368 17 2372
rect 21 2368 23 2372
rect 27 2368 29 2372
rect 33 2368 35 2372
rect 39 2368 41 2372
rect 45 2368 47 2372
rect 51 2368 53 2372
rect 57 2368 59 2372
rect 63 2368 65 2372
rect 69 2368 71 2372
rect 75 2368 77 2372
rect 81 2368 83 2372
rect 87 2368 89 2372
rect 93 2368 95 2372
rect 99 2368 101 2372
rect 105 2368 107 2372
rect 111 2368 113 2372
rect 117 2368 119 2372
rect 123 2368 125 2372
rect 129 2368 131 2372
rect 135 2368 137 2372
rect 141 2368 143 2372
rect 147 2368 149 2372
rect 153 2368 155 2372
rect 159 2368 161 2372
rect 165 2368 167 2372
rect 171 2368 173 2372
rect 177 2368 179 2372
rect 183 2368 185 2372
rect 189 2368 191 2372
rect 195 2368 197 2372
rect 201 2368 203 2372
rect 207 2368 209 2372
rect 213 2368 215 2372
rect 219 2368 221 2372
rect 225 2368 227 2372
rect 231 2368 233 2372
rect 237 2368 239 2372
rect 243 2368 245 2372
rect 249 2368 251 2372
rect 255 2368 257 2372
rect 261 2368 263 2372
rect 267 2368 269 2372
rect 273 2368 275 2372
rect 279 2368 281 2372
rect 285 2368 287 2372
rect 291 2368 293 2372
rect 297 2368 299 2372
rect 303 2368 305 2372
rect 309 2368 311 2372
rect 315 2368 317 2372
rect 321 2368 323 2372
rect 327 2368 329 2372
rect 333 2368 335 2372
rect 339 2368 341 2372
rect 345 2368 347 2372
rect 351 2368 353 2372
rect 357 2368 359 2372
rect 363 2368 365 2372
rect 365 2366 369 2368
rect 365 2360 369 2362
rect 365 2354 369 2356
rect 365 2348 369 2350
rect 365 2342 369 2344
rect 365 2336 369 2338
rect 365 2330 369 2332
rect 365 2324 369 2326
rect 365 2318 369 2320
rect 365 2312 369 2314
rect 365 2306 369 2308
rect 365 2300 369 2302
rect 365 2294 369 2296
rect 365 2288 369 2290
rect 365 2282 369 2284
rect 365 2276 369 2278
rect 365 2270 369 2272
rect 365 2264 369 2266
rect 365 2258 369 2260
rect 365 2252 369 2254
rect 365 2246 369 2248
rect 365 2240 372 2242
rect 369 2238 372 2240
rect 376 2238 412 2242
rect 421 2238 423 2242
rect 427 2238 429 2242
rect 433 2238 435 2242
rect 439 2238 441 2242
rect 450 2238 501 2242
rect 505 2238 509 2242
rect 369 2236 513 2238
rect 365 2234 372 2236
rect 369 2232 372 2234
rect 376 2232 412 2236
rect 421 2232 423 2236
rect 427 2232 429 2236
rect 433 2232 435 2236
rect 439 2232 441 2236
rect 450 2232 501 2236
rect 505 2232 509 2236
rect 369 2230 513 2232
rect 365 2228 372 2230
rect 369 2226 372 2228
rect 376 2226 412 2230
rect 421 2226 423 2230
rect 427 2226 429 2230
rect 433 2226 435 2230
rect 439 2226 441 2230
rect 450 2226 501 2230
rect 505 2226 509 2230
rect 369 2224 513 2226
rect 365 2222 372 2224
rect 369 2220 372 2222
rect 376 2220 412 2224
rect 421 2220 423 2224
rect 427 2220 429 2224
rect 433 2220 435 2224
rect 439 2220 441 2224
rect 450 2220 501 2224
rect 505 2220 509 2224
rect 369 2218 513 2220
rect 365 2216 372 2218
rect 369 2214 372 2216
rect 376 2214 412 2218
rect 421 2214 423 2218
rect 427 2214 429 2218
rect 433 2214 435 2218
rect 439 2214 441 2218
rect 450 2214 501 2218
rect 505 2214 509 2218
rect 369 2212 513 2214
rect 365 2210 372 2212
rect 369 2208 372 2210
rect 376 2208 412 2212
rect 421 2208 423 2212
rect 427 2208 429 2212
rect 433 2208 435 2212
rect 439 2208 441 2212
rect 450 2208 501 2212
rect 505 2208 509 2212
rect 369 2206 513 2208
rect 365 2204 372 2206
rect 369 2202 372 2204
rect 376 2202 412 2206
rect 421 2202 423 2206
rect 427 2202 429 2206
rect 433 2202 435 2206
rect 439 2202 441 2206
rect 450 2202 501 2206
rect 505 2202 509 2206
rect 365 2198 369 2200
rect 365 2192 369 2194
rect 388 2194 390 2198
rect 394 2194 397 2198
rect 401 2194 402 2198
rect 384 2192 406 2194
rect 365 2186 369 2188
rect 365 2180 369 2182
rect 365 2174 369 2176
rect 365 2168 369 2170
rect 365 2162 369 2164
rect 382 2188 384 2192
rect 388 2188 390 2192
rect 394 2188 397 2192
rect 401 2188 402 2192
rect 378 2186 406 2188
rect 382 2182 384 2186
rect 388 2182 390 2186
rect 394 2182 397 2186
rect 401 2182 402 2186
rect 378 2180 406 2182
rect 382 2176 384 2180
rect 388 2176 390 2180
rect 394 2176 397 2180
rect 401 2176 402 2180
rect 378 2174 406 2176
rect 382 2170 384 2174
rect 388 2170 390 2174
rect 394 2170 397 2174
rect 401 2170 402 2174
rect 378 2168 406 2170
rect 413 2197 465 2198
rect 413 2193 414 2197
rect 418 2193 420 2197
rect 424 2193 427 2197
rect 431 2193 433 2197
rect 437 2193 439 2197
rect 443 2193 445 2197
rect 449 2194 465 2197
rect 469 2194 471 2198
rect 475 2194 477 2198
rect 481 2194 483 2198
rect 487 2194 489 2198
rect 493 2194 509 2198
rect 449 2193 513 2194
rect 413 2192 513 2193
rect 413 2191 465 2192
rect 413 2187 414 2191
rect 418 2187 420 2191
rect 424 2187 427 2191
rect 431 2187 433 2191
rect 437 2187 439 2191
rect 443 2187 445 2191
rect 449 2188 465 2191
rect 469 2188 471 2192
rect 475 2188 477 2192
rect 481 2188 483 2192
rect 487 2188 489 2192
rect 493 2188 495 2192
rect 499 2188 509 2192
rect 449 2187 513 2188
rect 413 2186 513 2187
rect 413 2185 465 2186
rect 413 2181 414 2185
rect 418 2181 420 2185
rect 424 2181 427 2185
rect 431 2181 433 2185
rect 437 2181 439 2185
rect 443 2181 445 2185
rect 449 2182 465 2185
rect 469 2182 471 2186
rect 475 2182 477 2186
rect 481 2182 483 2186
rect 487 2182 489 2186
rect 493 2182 495 2186
rect 499 2182 509 2186
rect 449 2181 513 2182
rect 413 2180 513 2181
rect 413 2179 465 2180
rect 413 2175 414 2179
rect 418 2175 420 2179
rect 424 2175 427 2179
rect 431 2175 433 2179
rect 437 2175 439 2179
rect 443 2175 445 2179
rect 449 2176 465 2179
rect 469 2176 471 2180
rect 475 2176 477 2180
rect 481 2176 483 2180
rect 487 2176 489 2180
rect 493 2176 495 2180
rect 499 2176 509 2180
rect 449 2175 513 2176
rect 413 2174 513 2175
rect 413 2173 465 2174
rect 413 2169 414 2173
rect 418 2169 420 2173
rect 424 2169 427 2173
rect 431 2169 433 2173
rect 437 2169 439 2173
rect 443 2169 445 2173
rect 449 2170 465 2173
rect 469 2170 471 2174
rect 475 2170 477 2174
rect 481 2170 483 2174
rect 487 2170 489 2174
rect 493 2170 495 2174
rect 499 2170 509 2174
rect 449 2169 513 2170
rect 413 2168 513 2169
rect 382 2164 384 2168
rect 388 2164 390 2168
rect 394 2164 397 2168
rect 401 2164 402 2168
rect 469 2164 471 2168
rect 475 2164 477 2168
rect 481 2164 483 2168
rect 487 2164 489 2168
rect 493 2164 495 2168
rect 499 2164 509 2168
rect 378 2162 406 2164
rect 382 2158 384 2162
rect 388 2158 390 2162
rect 394 2158 397 2162
rect 401 2158 402 2162
rect 455 2160 456 2164
rect 460 2160 461 2164
rect 455 2159 461 2160
rect 365 2156 369 2158
rect 365 2150 369 2152
rect 455 2155 456 2159
rect 460 2155 461 2159
rect 465 2162 513 2164
rect 469 2158 471 2162
rect 475 2158 477 2162
rect 481 2158 483 2162
rect 487 2158 489 2162
rect 493 2158 495 2162
rect 499 2158 509 2162
rect 455 2154 461 2155
rect 455 2150 456 2154
rect 460 2150 509 2154
rect 455 2149 509 2150
rect 455 2145 456 2149
rect 460 2145 509 2149
rect 365 2114 369 2116
rect 365 2108 369 2110
rect 455 2117 456 2121
rect 460 2117 509 2121
rect 455 2116 509 2117
rect 455 2112 456 2116
rect 460 2112 509 2116
rect 455 2111 461 2112
rect 365 2102 369 2104
rect 365 2096 369 2098
rect 365 2090 369 2092
rect 365 2084 369 2086
rect 365 2078 369 2080
rect 382 2104 384 2108
rect 388 2104 390 2108
rect 394 2104 397 2108
rect 401 2104 402 2108
rect 378 2102 406 2104
rect 455 2107 456 2111
rect 460 2107 461 2111
rect 455 2106 461 2107
rect 455 2102 456 2106
rect 460 2102 461 2106
rect 469 2104 471 2108
rect 475 2104 477 2108
rect 481 2104 483 2108
rect 487 2104 489 2108
rect 493 2104 495 2108
rect 499 2104 509 2108
rect 465 2102 513 2104
rect 382 2098 384 2102
rect 388 2098 390 2102
rect 394 2098 397 2102
rect 401 2098 402 2102
rect 469 2098 471 2102
rect 475 2098 477 2102
rect 481 2098 483 2102
rect 487 2098 489 2102
rect 493 2098 495 2102
rect 499 2098 509 2102
rect 378 2096 406 2098
rect 382 2092 384 2096
rect 388 2092 390 2096
rect 394 2092 397 2096
rect 401 2092 402 2096
rect 378 2090 406 2092
rect 382 2086 384 2090
rect 388 2086 390 2090
rect 394 2086 397 2090
rect 401 2086 402 2090
rect 378 2084 406 2086
rect 382 2080 384 2084
rect 388 2080 390 2084
rect 394 2080 397 2084
rect 401 2080 402 2084
rect 378 2078 406 2080
rect 382 2074 384 2078
rect 388 2074 390 2078
rect 394 2074 397 2078
rect 401 2074 402 2078
rect 365 2072 369 2074
rect 384 2072 406 2074
rect 388 2068 390 2072
rect 394 2068 397 2072
rect 401 2068 402 2072
rect 413 2097 513 2098
rect 413 2093 414 2097
rect 418 2093 420 2097
rect 424 2093 427 2097
rect 431 2093 433 2097
rect 437 2093 439 2097
rect 443 2093 445 2097
rect 449 2096 513 2097
rect 449 2093 465 2096
rect 413 2092 465 2093
rect 469 2092 471 2096
rect 475 2092 477 2096
rect 481 2092 483 2096
rect 487 2092 489 2096
rect 493 2092 495 2096
rect 499 2092 509 2096
rect 413 2091 513 2092
rect 413 2087 414 2091
rect 418 2087 420 2091
rect 424 2087 427 2091
rect 431 2087 433 2091
rect 437 2087 439 2091
rect 443 2087 445 2091
rect 449 2090 513 2091
rect 449 2087 465 2090
rect 413 2086 465 2087
rect 469 2086 471 2090
rect 475 2086 477 2090
rect 481 2086 483 2090
rect 487 2086 489 2090
rect 493 2086 495 2090
rect 499 2086 509 2090
rect 413 2085 513 2086
rect 413 2081 414 2085
rect 418 2081 420 2085
rect 424 2081 427 2085
rect 431 2081 433 2085
rect 437 2081 439 2085
rect 443 2081 445 2085
rect 449 2084 513 2085
rect 449 2081 465 2084
rect 413 2080 465 2081
rect 469 2080 471 2084
rect 475 2080 477 2084
rect 481 2080 483 2084
rect 487 2080 489 2084
rect 493 2080 495 2084
rect 499 2080 509 2084
rect 413 2079 513 2080
rect 413 2075 414 2079
rect 418 2075 420 2079
rect 424 2075 427 2079
rect 431 2075 433 2079
rect 437 2075 439 2079
rect 443 2075 445 2079
rect 449 2078 513 2079
rect 449 2075 465 2078
rect 413 2074 465 2075
rect 469 2074 471 2078
rect 475 2074 477 2078
rect 481 2074 483 2078
rect 487 2074 489 2078
rect 493 2074 495 2078
rect 499 2074 509 2078
rect 413 2073 513 2074
rect 413 2069 414 2073
rect 418 2069 420 2073
rect 424 2069 427 2073
rect 431 2069 433 2073
rect 437 2069 439 2073
rect 443 2069 445 2073
rect 449 2072 513 2073
rect 449 2069 465 2072
rect 413 2068 465 2069
rect 469 2068 471 2072
rect 475 2068 477 2072
rect 481 2068 483 2072
rect 487 2068 489 2072
rect 493 2068 509 2072
rect 365 2066 369 2068
rect 369 2062 372 2064
rect 365 2060 372 2062
rect 376 2060 412 2064
rect 421 2060 423 2064
rect 427 2060 429 2064
rect 433 2060 435 2064
rect 439 2060 441 2064
rect 450 2060 501 2064
rect 505 2060 509 2064
rect 369 2058 513 2060
rect 369 2056 372 2058
rect 365 2054 372 2056
rect 376 2054 412 2058
rect 421 2054 423 2058
rect 427 2054 429 2058
rect 433 2054 435 2058
rect 439 2054 441 2058
rect 450 2054 501 2058
rect 505 2054 509 2058
rect 369 2052 513 2054
rect 369 2050 372 2052
rect 365 2048 372 2050
rect 376 2048 412 2052
rect 421 2048 423 2052
rect 427 2048 429 2052
rect 433 2048 435 2052
rect 439 2048 441 2052
rect 450 2048 501 2052
rect 505 2048 509 2052
rect 369 2046 513 2048
rect 369 2044 372 2046
rect 365 2042 372 2044
rect 376 2042 412 2046
rect 421 2042 423 2046
rect 427 2042 429 2046
rect 433 2042 435 2046
rect 439 2042 441 2046
rect 450 2042 501 2046
rect 505 2042 509 2046
rect 369 2040 513 2042
rect 369 2038 372 2040
rect 365 2036 372 2038
rect 376 2036 412 2040
rect 421 2036 423 2040
rect 427 2036 429 2040
rect 433 2036 435 2040
rect 439 2036 441 2040
rect 450 2036 501 2040
rect 505 2036 509 2040
rect 369 2034 513 2036
rect 369 2032 372 2034
rect 365 2030 372 2032
rect 376 2030 412 2034
rect 421 2030 423 2034
rect 427 2030 429 2034
rect 433 2030 435 2034
rect 439 2030 441 2034
rect 450 2030 501 2034
rect 505 2030 509 2034
rect 369 2028 513 2030
rect 369 2026 372 2028
rect 365 2024 372 2026
rect 376 2024 412 2028
rect 421 2024 423 2028
rect 427 2024 429 2028
rect 433 2024 435 2028
rect 439 2024 441 2028
rect 450 2024 501 2028
rect 505 2024 509 2028
rect 365 2018 369 2020
rect 365 2012 369 2014
rect 365 2006 369 2008
rect 365 2000 369 2002
rect 365 1994 369 1996
rect 365 1988 369 1990
rect 365 1982 369 1984
rect 365 1976 369 1978
rect 365 1970 369 1972
rect 365 1964 369 1966
rect 365 1958 369 1960
rect 365 1952 369 1954
rect 365 1946 369 1948
rect 365 1940 369 1942
rect 365 1934 369 1936
rect 365 1928 369 1930
rect 365 1922 369 1924
rect 365 1916 369 1918
rect 365 1910 369 1912
rect 365 1904 369 1906
rect 365 1898 369 1900
rect 3 1894 5 1898
rect 9 1894 11 1898
rect 15 1894 17 1898
rect 21 1894 23 1898
rect 27 1894 29 1898
rect 33 1894 35 1898
rect 39 1894 41 1898
rect 45 1894 47 1898
rect 51 1894 53 1898
rect 57 1894 59 1898
rect 63 1894 65 1898
rect 69 1894 71 1898
rect 75 1894 77 1898
rect 81 1894 83 1898
rect 87 1894 89 1898
rect 93 1894 95 1898
rect 99 1894 101 1898
rect 105 1894 107 1898
rect 111 1894 113 1898
rect 117 1894 119 1898
rect 123 1894 125 1898
rect 129 1894 131 1898
rect 135 1894 137 1898
rect 141 1894 143 1898
rect 147 1894 149 1898
rect 153 1894 155 1898
rect 159 1894 161 1898
rect 165 1894 167 1898
rect 171 1894 173 1898
rect 177 1894 179 1898
rect 183 1894 185 1898
rect 189 1894 191 1898
rect 195 1894 197 1898
rect 201 1894 203 1898
rect 207 1894 209 1898
rect 213 1894 215 1898
rect 219 1894 221 1898
rect 225 1894 227 1898
rect 231 1894 233 1898
rect 237 1894 239 1898
rect 243 1894 245 1898
rect 249 1894 251 1898
rect 255 1894 257 1898
rect 261 1894 263 1898
rect 267 1894 269 1898
rect 273 1894 275 1898
rect 279 1894 281 1898
rect 285 1894 287 1898
rect 291 1894 293 1898
rect 297 1894 299 1898
rect 303 1894 305 1898
rect 309 1894 311 1898
rect 315 1894 317 1898
rect 321 1894 323 1898
rect 327 1894 329 1898
rect 333 1894 335 1898
rect 339 1894 341 1898
rect 345 1894 347 1898
rect 351 1894 353 1898
rect 357 1894 359 1898
rect 363 1894 365 1898
rect 365 1892 369 1894
rect 365 1886 369 1888
rect 365 1880 369 1882
rect 365 1874 369 1876
rect 365 1868 369 1870
rect 365 1862 369 1864
rect 365 1856 369 1858
rect 365 1850 369 1852
rect 365 1844 369 1846
rect 365 1838 369 1840
rect 365 1832 369 1834
rect 365 1826 369 1828
rect 365 1820 369 1822
rect 365 1814 369 1816
rect 365 1808 369 1810
rect 365 1802 369 1804
rect 365 1796 369 1798
rect 365 1790 369 1792
rect 365 1784 369 1786
rect 365 1778 369 1780
rect 365 1772 369 1774
rect 365 1766 372 1768
rect 369 1764 372 1766
rect 376 1764 412 1768
rect 421 1764 423 1768
rect 427 1764 429 1768
rect 433 1764 435 1768
rect 439 1764 441 1768
rect 450 1764 501 1768
rect 505 1764 509 1768
rect 369 1762 513 1764
rect 365 1760 372 1762
rect 369 1758 372 1760
rect 376 1758 412 1762
rect 421 1758 423 1762
rect 427 1758 429 1762
rect 433 1758 435 1762
rect 439 1758 441 1762
rect 450 1758 501 1762
rect 505 1758 509 1762
rect 369 1756 513 1758
rect 365 1754 372 1756
rect 369 1752 372 1754
rect 376 1752 412 1756
rect 421 1752 423 1756
rect 427 1752 429 1756
rect 433 1752 435 1756
rect 439 1752 441 1756
rect 450 1752 501 1756
rect 505 1752 509 1756
rect 369 1750 513 1752
rect 365 1748 372 1750
rect 369 1746 372 1748
rect 376 1746 412 1750
rect 421 1746 423 1750
rect 427 1746 429 1750
rect 433 1746 435 1750
rect 439 1746 441 1750
rect 450 1746 501 1750
rect 505 1746 509 1750
rect 369 1744 513 1746
rect 365 1742 372 1744
rect 369 1740 372 1742
rect 376 1740 412 1744
rect 421 1740 423 1744
rect 427 1740 429 1744
rect 433 1740 435 1744
rect 439 1740 441 1744
rect 450 1740 501 1744
rect 505 1740 509 1744
rect 369 1738 513 1740
rect 365 1736 372 1738
rect 369 1734 372 1736
rect 376 1734 412 1738
rect 421 1734 423 1738
rect 427 1734 429 1738
rect 433 1734 435 1738
rect 439 1734 441 1738
rect 450 1734 501 1738
rect 505 1734 509 1738
rect 369 1732 513 1734
rect 365 1730 372 1732
rect 369 1728 372 1730
rect 376 1728 412 1732
rect 421 1728 423 1732
rect 427 1728 429 1732
rect 433 1728 435 1732
rect 439 1728 441 1732
rect 450 1728 501 1732
rect 505 1728 509 1732
rect 365 1724 369 1726
rect 365 1718 369 1720
rect 388 1720 390 1724
rect 394 1720 397 1724
rect 401 1720 402 1724
rect 384 1718 406 1720
rect 365 1712 369 1714
rect 365 1706 369 1708
rect 365 1700 369 1702
rect 365 1694 369 1696
rect 365 1688 369 1690
rect 382 1714 384 1718
rect 388 1714 390 1718
rect 394 1714 397 1718
rect 401 1714 402 1718
rect 378 1712 406 1714
rect 382 1708 384 1712
rect 388 1708 390 1712
rect 394 1708 397 1712
rect 401 1708 402 1712
rect 378 1706 406 1708
rect 382 1702 384 1706
rect 388 1702 390 1706
rect 394 1702 397 1706
rect 401 1702 402 1706
rect 378 1700 406 1702
rect 382 1696 384 1700
rect 388 1696 390 1700
rect 394 1696 397 1700
rect 401 1696 402 1700
rect 378 1694 406 1696
rect 413 1723 465 1724
rect 413 1719 414 1723
rect 418 1719 420 1723
rect 424 1719 427 1723
rect 431 1719 433 1723
rect 437 1719 439 1723
rect 443 1719 445 1723
rect 449 1720 465 1723
rect 469 1720 471 1724
rect 475 1720 477 1724
rect 481 1720 483 1724
rect 487 1720 489 1724
rect 493 1720 509 1724
rect 449 1719 513 1720
rect 413 1718 513 1719
rect 413 1717 465 1718
rect 413 1713 414 1717
rect 418 1713 420 1717
rect 424 1713 427 1717
rect 431 1713 433 1717
rect 437 1713 439 1717
rect 443 1713 445 1717
rect 449 1714 465 1717
rect 469 1714 471 1718
rect 475 1714 477 1718
rect 481 1714 483 1718
rect 487 1714 489 1718
rect 493 1714 495 1718
rect 499 1714 509 1718
rect 449 1713 513 1714
rect 413 1712 513 1713
rect 413 1711 465 1712
rect 413 1707 414 1711
rect 418 1707 420 1711
rect 424 1707 427 1711
rect 431 1707 433 1711
rect 437 1707 439 1711
rect 443 1707 445 1711
rect 449 1708 465 1711
rect 469 1708 471 1712
rect 475 1708 477 1712
rect 481 1708 483 1712
rect 487 1708 489 1712
rect 493 1708 495 1712
rect 499 1708 509 1712
rect 449 1707 513 1708
rect 413 1706 513 1707
rect 413 1705 465 1706
rect 413 1701 414 1705
rect 418 1701 420 1705
rect 424 1701 427 1705
rect 431 1701 433 1705
rect 437 1701 439 1705
rect 443 1701 445 1705
rect 449 1702 465 1705
rect 469 1702 471 1706
rect 475 1702 477 1706
rect 481 1702 483 1706
rect 487 1702 489 1706
rect 493 1702 495 1706
rect 499 1702 509 1706
rect 449 1701 513 1702
rect 413 1700 513 1701
rect 413 1699 465 1700
rect 413 1695 414 1699
rect 418 1695 420 1699
rect 424 1695 427 1699
rect 431 1695 433 1699
rect 437 1695 439 1699
rect 443 1695 445 1699
rect 449 1696 465 1699
rect 469 1696 471 1700
rect 475 1696 477 1700
rect 481 1696 483 1700
rect 487 1696 489 1700
rect 493 1696 495 1700
rect 499 1696 509 1700
rect 449 1695 513 1696
rect 413 1694 513 1695
rect 382 1690 384 1694
rect 388 1690 390 1694
rect 394 1690 397 1694
rect 401 1690 402 1694
rect 469 1690 471 1694
rect 475 1690 477 1694
rect 481 1690 483 1694
rect 487 1690 489 1694
rect 493 1690 495 1694
rect 499 1690 509 1694
rect 378 1688 406 1690
rect 382 1684 384 1688
rect 388 1684 390 1688
rect 394 1684 397 1688
rect 401 1684 402 1688
rect 455 1686 456 1690
rect 460 1686 461 1690
rect 455 1685 461 1686
rect 365 1682 369 1684
rect 365 1676 369 1678
rect 455 1681 456 1685
rect 460 1681 461 1685
rect 465 1688 513 1690
rect 469 1684 471 1688
rect 475 1684 477 1688
rect 481 1684 483 1688
rect 487 1684 489 1688
rect 493 1684 495 1688
rect 499 1684 509 1688
rect 455 1680 461 1681
rect 455 1676 456 1680
rect 460 1676 509 1680
rect 455 1675 509 1676
rect 455 1671 456 1675
rect 460 1671 509 1675
rect 365 1640 369 1642
rect 365 1634 369 1636
rect 455 1643 456 1647
rect 460 1643 509 1647
rect 455 1642 509 1643
rect 455 1638 456 1642
rect 460 1638 509 1642
rect 455 1637 461 1638
rect 365 1628 369 1630
rect 365 1622 369 1624
rect 365 1616 369 1618
rect 365 1610 369 1612
rect 365 1604 369 1606
rect 382 1630 384 1634
rect 388 1630 390 1634
rect 394 1630 397 1634
rect 401 1630 402 1634
rect 378 1628 406 1630
rect 455 1633 456 1637
rect 460 1633 461 1637
rect 455 1632 461 1633
rect 455 1628 456 1632
rect 460 1628 461 1632
rect 469 1630 471 1634
rect 475 1630 477 1634
rect 481 1630 483 1634
rect 487 1630 489 1634
rect 493 1630 495 1634
rect 499 1630 509 1634
rect 465 1628 513 1630
rect 382 1624 384 1628
rect 388 1624 390 1628
rect 394 1624 397 1628
rect 401 1624 402 1628
rect 469 1624 471 1628
rect 475 1624 477 1628
rect 481 1624 483 1628
rect 487 1624 489 1628
rect 493 1624 495 1628
rect 499 1624 509 1628
rect 378 1622 406 1624
rect 382 1618 384 1622
rect 388 1618 390 1622
rect 394 1618 397 1622
rect 401 1618 402 1622
rect 378 1616 406 1618
rect 382 1612 384 1616
rect 388 1612 390 1616
rect 394 1612 397 1616
rect 401 1612 402 1616
rect 378 1610 406 1612
rect 382 1606 384 1610
rect 388 1606 390 1610
rect 394 1606 397 1610
rect 401 1606 402 1610
rect 378 1604 406 1606
rect 382 1600 384 1604
rect 388 1600 390 1604
rect 394 1600 397 1604
rect 401 1600 402 1604
rect 365 1598 369 1600
rect 384 1598 406 1600
rect 388 1594 390 1598
rect 394 1594 397 1598
rect 401 1594 402 1598
rect 413 1623 513 1624
rect 413 1619 414 1623
rect 418 1619 420 1623
rect 424 1619 427 1623
rect 431 1619 433 1623
rect 437 1619 439 1623
rect 443 1619 445 1623
rect 449 1622 513 1623
rect 449 1619 465 1622
rect 413 1618 465 1619
rect 469 1618 471 1622
rect 475 1618 477 1622
rect 481 1618 483 1622
rect 487 1618 489 1622
rect 493 1618 495 1622
rect 499 1618 509 1622
rect 413 1617 513 1618
rect 413 1613 414 1617
rect 418 1613 420 1617
rect 424 1613 427 1617
rect 431 1613 433 1617
rect 437 1613 439 1617
rect 443 1613 445 1617
rect 449 1616 513 1617
rect 449 1613 465 1616
rect 413 1612 465 1613
rect 469 1612 471 1616
rect 475 1612 477 1616
rect 481 1612 483 1616
rect 487 1612 489 1616
rect 493 1612 495 1616
rect 499 1612 509 1616
rect 413 1611 513 1612
rect 413 1607 414 1611
rect 418 1607 420 1611
rect 424 1607 427 1611
rect 431 1607 433 1611
rect 437 1607 439 1611
rect 443 1607 445 1611
rect 449 1610 513 1611
rect 449 1607 465 1610
rect 413 1606 465 1607
rect 469 1606 471 1610
rect 475 1606 477 1610
rect 481 1606 483 1610
rect 487 1606 489 1610
rect 493 1606 495 1610
rect 499 1606 509 1610
rect 413 1605 513 1606
rect 413 1601 414 1605
rect 418 1601 420 1605
rect 424 1601 427 1605
rect 431 1601 433 1605
rect 437 1601 439 1605
rect 443 1601 445 1605
rect 449 1604 513 1605
rect 449 1601 465 1604
rect 413 1600 465 1601
rect 469 1600 471 1604
rect 475 1600 477 1604
rect 481 1600 483 1604
rect 487 1600 489 1604
rect 493 1600 495 1604
rect 499 1600 509 1604
rect 413 1599 513 1600
rect 413 1595 414 1599
rect 418 1595 420 1599
rect 424 1595 427 1599
rect 431 1595 433 1599
rect 437 1595 439 1599
rect 443 1595 445 1599
rect 449 1598 513 1599
rect 449 1595 465 1598
rect 413 1594 465 1595
rect 469 1594 471 1598
rect 475 1594 477 1598
rect 481 1594 483 1598
rect 487 1594 489 1598
rect 493 1594 509 1598
rect 365 1592 369 1594
rect 369 1588 372 1590
rect 365 1586 372 1588
rect 376 1586 412 1590
rect 421 1586 423 1590
rect 427 1586 429 1590
rect 433 1586 435 1590
rect 439 1586 441 1590
rect 450 1586 501 1590
rect 505 1586 509 1590
rect 369 1584 513 1586
rect 369 1582 372 1584
rect 365 1580 372 1582
rect 376 1580 412 1584
rect 421 1580 423 1584
rect 427 1580 429 1584
rect 433 1580 435 1584
rect 439 1580 441 1584
rect 450 1580 501 1584
rect 505 1580 509 1584
rect 369 1578 513 1580
rect 369 1576 372 1578
rect 365 1574 372 1576
rect 376 1574 412 1578
rect 421 1574 423 1578
rect 427 1574 429 1578
rect 433 1574 435 1578
rect 439 1574 441 1578
rect 450 1574 501 1578
rect 505 1574 509 1578
rect 369 1572 513 1574
rect 369 1570 372 1572
rect 365 1568 372 1570
rect 376 1568 412 1572
rect 421 1568 423 1572
rect 427 1568 429 1572
rect 433 1568 435 1572
rect 439 1568 441 1572
rect 450 1568 501 1572
rect 505 1568 509 1572
rect 369 1566 513 1568
rect 369 1564 372 1566
rect 365 1562 372 1564
rect 376 1562 412 1566
rect 421 1562 423 1566
rect 427 1562 429 1566
rect 433 1562 435 1566
rect 439 1562 441 1566
rect 450 1562 501 1566
rect 505 1562 509 1566
rect 369 1560 513 1562
rect 369 1558 372 1560
rect 365 1556 372 1558
rect 376 1556 412 1560
rect 421 1556 423 1560
rect 427 1556 429 1560
rect 433 1556 435 1560
rect 439 1556 441 1560
rect 450 1556 501 1560
rect 505 1556 509 1560
rect 369 1554 513 1556
rect 369 1552 372 1554
rect 365 1550 372 1552
rect 376 1550 412 1554
rect 421 1550 423 1554
rect 427 1550 429 1554
rect 433 1550 435 1554
rect 439 1550 441 1554
rect 450 1550 501 1554
rect 505 1550 509 1554
rect 365 1544 369 1546
rect 365 1538 369 1540
rect 365 1532 369 1534
rect 365 1526 369 1528
rect 365 1520 369 1522
rect 365 1514 369 1516
rect 365 1508 369 1510
rect 365 1502 369 1504
rect 365 1496 369 1498
rect 365 1490 369 1492
rect 365 1484 369 1486
rect 365 1478 369 1480
rect 365 1472 369 1474
rect 365 1466 369 1468
rect 365 1460 369 1462
rect 365 1454 369 1456
rect 365 1448 369 1450
rect 365 1442 369 1444
rect 365 1436 369 1438
rect 365 1430 369 1432
rect 365 1424 369 1426
rect 3 1420 5 1424
rect 9 1420 11 1424
rect 15 1420 17 1424
rect 21 1420 23 1424
rect 27 1420 29 1424
rect 33 1420 35 1424
rect 39 1420 41 1424
rect 45 1420 47 1424
rect 51 1420 53 1424
rect 57 1420 59 1424
rect 63 1420 65 1424
rect 69 1420 71 1424
rect 75 1420 77 1424
rect 81 1420 83 1424
rect 87 1420 89 1424
rect 93 1420 95 1424
rect 99 1420 101 1424
rect 105 1420 107 1424
rect 111 1420 113 1424
rect 117 1420 119 1424
rect 123 1420 125 1424
rect 129 1420 131 1424
rect 135 1420 137 1424
rect 141 1420 143 1424
rect 147 1420 149 1424
rect 153 1420 155 1424
rect 159 1420 161 1424
rect 165 1420 167 1424
rect 171 1420 173 1424
rect 177 1420 179 1424
rect 183 1420 185 1424
rect 189 1420 191 1424
rect 195 1420 197 1424
rect 201 1420 203 1424
rect 207 1420 209 1424
rect 213 1420 215 1424
rect 219 1420 221 1424
rect 225 1420 227 1424
rect 231 1420 233 1424
rect 237 1420 239 1424
rect 243 1420 245 1424
rect 249 1420 251 1424
rect 255 1420 257 1424
rect 261 1420 263 1424
rect 267 1420 269 1424
rect 273 1420 275 1424
rect 279 1420 281 1424
rect 285 1420 287 1424
rect 291 1420 293 1424
rect 297 1420 299 1424
rect 303 1420 305 1424
rect 309 1420 311 1424
rect 315 1420 317 1424
rect 321 1420 323 1424
rect 327 1420 329 1424
rect 333 1420 335 1424
rect 339 1420 341 1424
rect 345 1420 347 1424
rect 351 1420 353 1424
rect 357 1420 359 1424
rect 363 1420 365 1424
rect 365 1418 369 1420
rect 365 1412 369 1414
rect 365 1406 369 1408
rect 365 1400 369 1402
rect 365 1394 369 1396
rect 365 1388 369 1390
rect 365 1382 369 1384
rect 365 1376 369 1378
rect 365 1370 369 1372
rect 365 1364 369 1366
rect 365 1358 369 1360
rect 365 1352 369 1354
rect 365 1346 369 1348
rect 365 1340 369 1342
rect 365 1334 369 1336
rect 365 1328 369 1330
rect 365 1322 369 1324
rect 365 1316 369 1318
rect 365 1310 369 1312
rect 365 1304 369 1306
rect 365 1298 369 1300
rect 365 1292 372 1294
rect 369 1290 372 1292
rect 376 1290 412 1294
rect 421 1290 423 1294
rect 427 1290 429 1294
rect 433 1290 435 1294
rect 439 1290 441 1294
rect 450 1290 501 1294
rect 505 1290 509 1294
rect 369 1288 513 1290
rect 365 1286 372 1288
rect 369 1284 372 1286
rect 376 1284 412 1288
rect 421 1284 423 1288
rect 427 1284 429 1288
rect 433 1284 435 1288
rect 439 1284 441 1288
rect 450 1284 501 1288
rect 505 1284 509 1288
rect 369 1282 513 1284
rect 365 1280 372 1282
rect 369 1278 372 1280
rect 376 1278 412 1282
rect 421 1278 423 1282
rect 427 1278 429 1282
rect 433 1278 435 1282
rect 439 1278 441 1282
rect 450 1278 501 1282
rect 505 1278 509 1282
rect 369 1276 513 1278
rect 365 1274 372 1276
rect 369 1272 372 1274
rect 376 1272 412 1276
rect 421 1272 423 1276
rect 427 1272 429 1276
rect 433 1272 435 1276
rect 439 1272 441 1276
rect 450 1272 501 1276
rect 505 1272 509 1276
rect 369 1270 513 1272
rect 365 1268 372 1270
rect 369 1266 372 1268
rect 376 1266 412 1270
rect 421 1266 423 1270
rect 427 1266 429 1270
rect 433 1266 435 1270
rect 439 1266 441 1270
rect 450 1266 501 1270
rect 505 1266 509 1270
rect 369 1264 513 1266
rect 365 1262 372 1264
rect 369 1260 372 1262
rect 376 1260 412 1264
rect 421 1260 423 1264
rect 427 1260 429 1264
rect 433 1260 435 1264
rect 439 1260 441 1264
rect 450 1260 501 1264
rect 505 1260 509 1264
rect 369 1258 513 1260
rect 365 1256 372 1258
rect 369 1254 372 1256
rect 376 1254 412 1258
rect 421 1254 423 1258
rect 427 1254 429 1258
rect 433 1254 435 1258
rect 439 1254 441 1258
rect 450 1254 501 1258
rect 505 1254 509 1258
rect 365 1250 369 1252
rect 365 1244 369 1246
rect 388 1246 390 1250
rect 394 1246 397 1250
rect 401 1246 402 1250
rect 384 1244 406 1246
rect 365 1238 369 1240
rect 365 1232 369 1234
rect 365 1226 369 1228
rect 365 1220 369 1222
rect 365 1214 369 1216
rect 382 1240 384 1244
rect 388 1240 390 1244
rect 394 1240 397 1244
rect 401 1240 402 1244
rect 378 1238 406 1240
rect 382 1234 384 1238
rect 388 1234 390 1238
rect 394 1234 397 1238
rect 401 1234 402 1238
rect 378 1232 406 1234
rect 382 1228 384 1232
rect 388 1228 390 1232
rect 394 1228 397 1232
rect 401 1228 402 1232
rect 378 1226 406 1228
rect 382 1222 384 1226
rect 388 1222 390 1226
rect 394 1222 397 1226
rect 401 1222 402 1226
rect 378 1220 406 1222
rect 413 1249 465 1250
rect 413 1245 414 1249
rect 418 1245 420 1249
rect 424 1245 427 1249
rect 431 1245 433 1249
rect 437 1245 439 1249
rect 443 1245 445 1249
rect 449 1246 465 1249
rect 469 1246 471 1250
rect 475 1246 477 1250
rect 481 1246 483 1250
rect 487 1246 489 1250
rect 493 1246 509 1250
rect 449 1245 513 1246
rect 413 1244 513 1245
rect 413 1243 465 1244
rect 413 1239 414 1243
rect 418 1239 420 1243
rect 424 1239 427 1243
rect 431 1239 433 1243
rect 437 1239 439 1243
rect 443 1239 445 1243
rect 449 1240 465 1243
rect 469 1240 471 1244
rect 475 1240 477 1244
rect 481 1240 483 1244
rect 487 1240 489 1244
rect 493 1240 495 1244
rect 499 1240 509 1244
rect 449 1239 513 1240
rect 413 1238 513 1239
rect 413 1237 465 1238
rect 413 1233 414 1237
rect 418 1233 420 1237
rect 424 1233 427 1237
rect 431 1233 433 1237
rect 437 1233 439 1237
rect 443 1233 445 1237
rect 449 1234 465 1237
rect 469 1234 471 1238
rect 475 1234 477 1238
rect 481 1234 483 1238
rect 487 1234 489 1238
rect 493 1234 495 1238
rect 499 1234 509 1238
rect 449 1233 513 1234
rect 413 1232 513 1233
rect 413 1231 465 1232
rect 413 1227 414 1231
rect 418 1227 420 1231
rect 424 1227 427 1231
rect 431 1227 433 1231
rect 437 1227 439 1231
rect 443 1227 445 1231
rect 449 1228 465 1231
rect 469 1228 471 1232
rect 475 1228 477 1232
rect 481 1228 483 1232
rect 487 1228 489 1232
rect 493 1228 495 1232
rect 499 1228 509 1232
rect 449 1227 513 1228
rect 413 1226 513 1227
rect 413 1225 465 1226
rect 413 1221 414 1225
rect 418 1221 420 1225
rect 424 1221 427 1225
rect 431 1221 433 1225
rect 437 1221 439 1225
rect 443 1221 445 1225
rect 449 1222 465 1225
rect 469 1222 471 1226
rect 475 1222 477 1226
rect 481 1222 483 1226
rect 487 1222 489 1226
rect 493 1222 495 1226
rect 499 1222 509 1226
rect 449 1221 513 1222
rect 413 1220 513 1221
rect 382 1216 384 1220
rect 388 1216 390 1220
rect 394 1216 397 1220
rect 401 1216 402 1220
rect 469 1216 471 1220
rect 475 1216 477 1220
rect 481 1216 483 1220
rect 487 1216 489 1220
rect 493 1216 495 1220
rect 499 1216 509 1220
rect 378 1214 406 1216
rect 382 1210 384 1214
rect 388 1210 390 1214
rect 394 1210 397 1214
rect 401 1210 402 1214
rect 455 1212 456 1216
rect 460 1212 461 1216
rect 455 1211 461 1212
rect 365 1208 369 1210
rect 365 1202 369 1204
rect 455 1207 456 1211
rect 460 1207 461 1211
rect 465 1214 513 1216
rect 469 1210 471 1214
rect 475 1210 477 1214
rect 481 1210 483 1214
rect 487 1210 489 1214
rect 493 1210 495 1214
rect 499 1210 509 1214
rect 455 1206 461 1207
rect 455 1202 456 1206
rect 460 1202 509 1206
rect 455 1201 509 1202
rect 455 1197 456 1201
rect 460 1197 509 1201
rect 365 1166 369 1168
rect 365 1160 369 1162
rect 455 1169 456 1173
rect 460 1169 509 1173
rect 455 1168 509 1169
rect 455 1164 456 1168
rect 460 1164 509 1168
rect 455 1163 461 1164
rect 365 1154 369 1156
rect 365 1148 369 1150
rect 365 1142 369 1144
rect 365 1136 369 1138
rect 365 1130 369 1132
rect 382 1156 384 1160
rect 388 1156 390 1160
rect 394 1156 397 1160
rect 401 1156 402 1160
rect 378 1154 406 1156
rect 455 1159 456 1163
rect 460 1159 461 1163
rect 455 1158 461 1159
rect 455 1154 456 1158
rect 460 1154 461 1158
rect 469 1156 471 1160
rect 475 1156 477 1160
rect 481 1156 483 1160
rect 487 1156 489 1160
rect 493 1156 495 1160
rect 499 1156 509 1160
rect 465 1154 513 1156
rect 382 1150 384 1154
rect 388 1150 390 1154
rect 394 1150 397 1154
rect 401 1150 402 1154
rect 469 1150 471 1154
rect 475 1150 477 1154
rect 481 1150 483 1154
rect 487 1150 489 1154
rect 493 1150 495 1154
rect 499 1150 509 1154
rect 378 1148 406 1150
rect 382 1144 384 1148
rect 388 1144 390 1148
rect 394 1144 397 1148
rect 401 1144 402 1148
rect 378 1142 406 1144
rect 382 1138 384 1142
rect 388 1138 390 1142
rect 394 1138 397 1142
rect 401 1138 402 1142
rect 378 1136 406 1138
rect 382 1132 384 1136
rect 388 1132 390 1136
rect 394 1132 397 1136
rect 401 1132 402 1136
rect 378 1130 406 1132
rect 382 1126 384 1130
rect 388 1126 390 1130
rect 394 1126 397 1130
rect 401 1126 402 1130
rect 365 1124 369 1126
rect 384 1124 406 1126
rect 388 1120 390 1124
rect 394 1120 397 1124
rect 401 1120 402 1124
rect 413 1149 513 1150
rect 413 1145 414 1149
rect 418 1145 420 1149
rect 424 1145 427 1149
rect 431 1145 433 1149
rect 437 1145 439 1149
rect 443 1145 445 1149
rect 449 1148 513 1149
rect 449 1145 465 1148
rect 413 1144 465 1145
rect 469 1144 471 1148
rect 475 1144 477 1148
rect 481 1144 483 1148
rect 487 1144 489 1148
rect 493 1144 495 1148
rect 499 1144 509 1148
rect 413 1143 513 1144
rect 413 1139 414 1143
rect 418 1139 420 1143
rect 424 1139 427 1143
rect 431 1139 433 1143
rect 437 1139 439 1143
rect 443 1139 445 1143
rect 449 1142 513 1143
rect 449 1139 465 1142
rect 413 1138 465 1139
rect 469 1138 471 1142
rect 475 1138 477 1142
rect 481 1138 483 1142
rect 487 1138 489 1142
rect 493 1138 495 1142
rect 499 1138 509 1142
rect 413 1137 513 1138
rect 413 1133 414 1137
rect 418 1133 420 1137
rect 424 1133 427 1137
rect 431 1133 433 1137
rect 437 1133 439 1137
rect 443 1133 445 1137
rect 449 1136 513 1137
rect 449 1133 465 1136
rect 413 1132 465 1133
rect 469 1132 471 1136
rect 475 1132 477 1136
rect 481 1132 483 1136
rect 487 1132 489 1136
rect 493 1132 495 1136
rect 499 1132 509 1136
rect 413 1131 513 1132
rect 413 1127 414 1131
rect 418 1127 420 1131
rect 424 1127 427 1131
rect 431 1127 433 1131
rect 437 1127 439 1131
rect 443 1127 445 1131
rect 449 1130 513 1131
rect 449 1127 465 1130
rect 413 1126 465 1127
rect 469 1126 471 1130
rect 475 1126 477 1130
rect 481 1126 483 1130
rect 487 1126 489 1130
rect 493 1126 495 1130
rect 499 1126 509 1130
rect 413 1125 513 1126
rect 413 1121 414 1125
rect 418 1121 420 1125
rect 424 1121 427 1125
rect 431 1121 433 1125
rect 437 1121 439 1125
rect 443 1121 445 1125
rect 449 1124 513 1125
rect 449 1121 465 1124
rect 413 1120 465 1121
rect 469 1120 471 1124
rect 475 1120 477 1124
rect 481 1120 483 1124
rect 487 1120 489 1124
rect 493 1120 509 1124
rect 365 1118 369 1120
rect 369 1114 372 1116
rect 365 1112 372 1114
rect 376 1112 412 1116
rect 421 1112 423 1116
rect 427 1112 429 1116
rect 433 1112 435 1116
rect 439 1112 441 1116
rect 450 1112 501 1116
rect 505 1112 509 1116
rect 369 1110 513 1112
rect 369 1108 372 1110
rect 365 1106 372 1108
rect 376 1106 412 1110
rect 421 1106 423 1110
rect 427 1106 429 1110
rect 433 1106 435 1110
rect 439 1106 441 1110
rect 450 1106 501 1110
rect 505 1106 509 1110
rect 369 1104 513 1106
rect 369 1102 372 1104
rect 365 1100 372 1102
rect 376 1100 412 1104
rect 421 1100 423 1104
rect 427 1100 429 1104
rect 433 1100 435 1104
rect 439 1100 441 1104
rect 450 1100 501 1104
rect 505 1100 509 1104
rect 369 1098 513 1100
rect 369 1096 372 1098
rect 365 1094 372 1096
rect 376 1094 412 1098
rect 421 1094 423 1098
rect 427 1094 429 1098
rect 433 1094 435 1098
rect 439 1094 441 1098
rect 450 1094 501 1098
rect 505 1094 509 1098
rect 369 1092 513 1094
rect 369 1090 372 1092
rect 365 1088 372 1090
rect 376 1088 412 1092
rect 421 1088 423 1092
rect 427 1088 429 1092
rect 433 1088 435 1092
rect 439 1088 441 1092
rect 450 1088 501 1092
rect 505 1088 509 1092
rect 369 1086 513 1088
rect 369 1084 372 1086
rect 365 1082 372 1084
rect 376 1082 412 1086
rect 421 1082 423 1086
rect 427 1082 429 1086
rect 433 1082 435 1086
rect 439 1082 441 1086
rect 450 1082 501 1086
rect 505 1082 509 1086
rect 369 1080 513 1082
rect 369 1078 372 1080
rect 365 1076 372 1078
rect 376 1076 412 1080
rect 421 1076 423 1080
rect 427 1076 429 1080
rect 433 1076 435 1080
rect 439 1076 441 1080
rect 450 1076 501 1080
rect 505 1076 509 1080
rect 365 1070 369 1072
rect 365 1064 369 1066
rect 365 1058 369 1060
rect 365 1052 369 1054
rect 365 1046 369 1048
rect 365 1040 369 1042
rect 365 1034 369 1036
rect 365 1028 369 1030
rect 365 1022 369 1024
rect 365 1016 369 1018
rect 365 1010 369 1012
rect 365 1004 369 1006
rect 365 998 369 1000
rect 365 992 369 994
rect 365 986 369 988
rect 365 980 369 982
rect 365 974 369 976
rect 365 968 369 970
rect 365 962 369 964
rect 365 956 369 958
rect 365 950 369 952
rect 3 946 5 950
rect 9 946 11 950
rect 15 946 17 950
rect 21 946 23 950
rect 27 946 29 950
rect 33 946 35 950
rect 39 946 41 950
rect 45 946 47 950
rect 51 946 53 950
rect 57 946 59 950
rect 63 946 65 950
rect 69 946 71 950
rect 75 946 77 950
rect 81 946 83 950
rect 87 946 89 950
rect 93 946 95 950
rect 99 946 101 950
rect 105 946 107 950
rect 111 946 113 950
rect 117 946 119 950
rect 123 946 125 950
rect 129 946 131 950
rect 135 946 137 950
rect 141 946 143 950
rect 147 946 149 950
rect 153 946 155 950
rect 159 946 161 950
rect 165 946 167 950
rect 171 946 173 950
rect 177 946 179 950
rect 183 946 185 950
rect 189 946 191 950
rect 195 946 197 950
rect 201 946 203 950
rect 207 946 209 950
rect 213 946 215 950
rect 219 946 221 950
rect 225 946 227 950
rect 231 946 233 950
rect 237 946 239 950
rect 243 946 245 950
rect 249 946 251 950
rect 255 946 257 950
rect 261 946 263 950
rect 267 946 269 950
rect 273 946 275 950
rect 279 946 281 950
rect 285 946 287 950
rect 291 946 293 950
rect 297 946 299 950
rect 303 946 305 950
rect 309 946 311 950
rect 315 946 317 950
rect 321 946 323 950
rect 327 946 329 950
rect 333 946 335 950
rect 339 946 341 950
rect 345 946 347 950
rect 351 946 353 950
rect 357 946 359 950
rect 363 946 365 950
rect 365 944 369 946
rect 365 938 369 940
rect 365 932 369 934
rect 365 926 369 928
rect 365 920 369 922
rect 365 914 369 916
rect 365 908 369 910
rect 365 902 369 904
rect 365 896 369 898
rect 365 890 369 892
rect 365 884 369 886
rect 365 878 369 880
rect 365 872 369 874
rect 365 866 369 868
rect 365 860 369 862
rect 365 854 369 856
rect 365 848 369 850
rect 365 842 369 844
rect 365 836 369 838
rect 365 830 369 832
rect 365 824 369 826
rect 365 818 372 820
rect 369 816 372 818
rect 376 816 412 820
rect 421 816 423 820
rect 427 816 429 820
rect 433 816 435 820
rect 439 816 441 820
rect 450 816 501 820
rect 505 816 509 820
rect 369 814 513 816
rect 365 812 372 814
rect 369 810 372 812
rect 376 810 412 814
rect 421 810 423 814
rect 427 810 429 814
rect 433 810 435 814
rect 439 810 441 814
rect 450 810 501 814
rect 505 810 509 814
rect 369 808 513 810
rect 365 806 372 808
rect 369 804 372 806
rect 376 804 412 808
rect 421 804 423 808
rect 427 804 429 808
rect 433 804 435 808
rect 439 804 441 808
rect 450 804 501 808
rect 505 804 509 808
rect 369 802 513 804
rect 365 800 372 802
rect 369 798 372 800
rect 376 798 412 802
rect 421 798 423 802
rect 427 798 429 802
rect 433 798 435 802
rect 439 798 441 802
rect 450 798 501 802
rect 505 798 509 802
rect 369 796 513 798
rect 365 794 372 796
rect 369 792 372 794
rect 376 792 412 796
rect 421 792 423 796
rect 427 792 429 796
rect 433 792 435 796
rect 439 792 441 796
rect 450 792 501 796
rect 505 792 509 796
rect 369 790 513 792
rect 365 788 372 790
rect 369 786 372 788
rect 376 786 412 790
rect 421 786 423 790
rect 427 786 429 790
rect 433 786 435 790
rect 439 786 441 790
rect 450 786 501 790
rect 505 786 509 790
rect 369 784 513 786
rect 365 782 372 784
rect 369 780 372 782
rect 376 780 412 784
rect 421 780 423 784
rect 427 780 429 784
rect 433 780 435 784
rect 439 780 441 784
rect 450 780 501 784
rect 505 780 509 784
rect 365 776 369 778
rect 365 770 369 772
rect 388 772 390 776
rect 394 772 397 776
rect 401 772 402 776
rect 384 770 406 772
rect 365 764 369 766
rect 365 758 369 760
rect 365 752 369 754
rect 365 746 369 748
rect 365 740 369 742
rect 382 766 384 770
rect 388 766 390 770
rect 394 766 397 770
rect 401 766 402 770
rect 378 764 406 766
rect 382 760 384 764
rect 388 760 390 764
rect 394 760 397 764
rect 401 760 402 764
rect 378 758 406 760
rect 382 754 384 758
rect 388 754 390 758
rect 394 754 397 758
rect 401 754 402 758
rect 378 752 406 754
rect 382 748 384 752
rect 388 748 390 752
rect 394 748 397 752
rect 401 748 402 752
rect 378 746 406 748
rect 413 775 465 776
rect 413 771 414 775
rect 418 771 420 775
rect 424 771 427 775
rect 431 771 433 775
rect 437 771 439 775
rect 443 771 445 775
rect 449 772 465 775
rect 469 772 471 776
rect 475 772 477 776
rect 481 772 483 776
rect 487 772 489 776
rect 493 772 509 776
rect 449 771 513 772
rect 413 770 513 771
rect 413 769 465 770
rect 413 765 414 769
rect 418 765 420 769
rect 424 765 427 769
rect 431 765 433 769
rect 437 765 439 769
rect 443 765 445 769
rect 449 766 465 769
rect 469 766 471 770
rect 475 766 477 770
rect 481 766 483 770
rect 487 766 489 770
rect 493 766 495 770
rect 499 766 509 770
rect 449 765 513 766
rect 413 764 513 765
rect 413 763 465 764
rect 413 759 414 763
rect 418 759 420 763
rect 424 759 427 763
rect 431 759 433 763
rect 437 759 439 763
rect 443 759 445 763
rect 449 760 465 763
rect 469 760 471 764
rect 475 760 477 764
rect 481 760 483 764
rect 487 760 489 764
rect 493 760 495 764
rect 499 760 509 764
rect 449 759 513 760
rect 413 758 513 759
rect 413 757 465 758
rect 413 753 414 757
rect 418 753 420 757
rect 424 753 427 757
rect 431 753 433 757
rect 437 753 439 757
rect 443 753 445 757
rect 449 754 465 757
rect 469 754 471 758
rect 475 754 477 758
rect 481 754 483 758
rect 487 754 489 758
rect 493 754 495 758
rect 499 754 509 758
rect 449 753 513 754
rect 413 752 513 753
rect 413 751 465 752
rect 413 747 414 751
rect 418 747 420 751
rect 424 747 427 751
rect 431 747 433 751
rect 437 747 439 751
rect 443 747 445 751
rect 449 748 465 751
rect 469 748 471 752
rect 475 748 477 752
rect 481 748 483 752
rect 487 748 489 752
rect 493 748 495 752
rect 499 748 509 752
rect 449 747 513 748
rect 413 746 513 747
rect 382 742 384 746
rect 388 742 390 746
rect 394 742 397 746
rect 401 742 402 746
rect 469 742 471 746
rect 475 742 477 746
rect 481 742 483 746
rect 487 742 489 746
rect 493 742 495 746
rect 499 742 509 746
rect 378 740 406 742
rect 382 736 384 740
rect 388 736 390 740
rect 394 736 397 740
rect 401 736 402 740
rect 455 738 456 742
rect 460 738 461 742
rect 455 737 461 738
rect 365 734 369 736
rect 365 728 369 730
rect 455 733 456 737
rect 460 733 461 737
rect 465 740 513 742
rect 469 736 471 740
rect 475 736 477 740
rect 481 736 483 740
rect 487 736 489 740
rect 493 736 495 740
rect 499 736 509 740
rect 455 732 461 733
rect 455 728 456 732
rect 460 728 509 732
rect 455 727 509 728
rect 455 723 456 727
rect 460 723 509 727
rect 365 692 369 694
rect 365 686 369 688
rect 455 695 456 699
rect 460 695 509 699
rect 455 694 509 695
rect 455 690 456 694
rect 460 690 509 694
rect 455 689 461 690
rect 365 680 369 682
rect 365 674 369 676
rect 365 668 369 670
rect 365 662 369 664
rect 365 656 369 658
rect 382 682 384 686
rect 388 682 390 686
rect 394 682 397 686
rect 401 682 402 686
rect 378 680 406 682
rect 455 685 456 689
rect 460 685 461 689
rect 455 684 461 685
rect 455 680 456 684
rect 460 680 461 684
rect 469 682 471 686
rect 475 682 477 686
rect 481 682 483 686
rect 487 682 489 686
rect 493 682 495 686
rect 499 682 509 686
rect 465 680 513 682
rect 382 676 384 680
rect 388 676 390 680
rect 394 676 397 680
rect 401 676 402 680
rect 469 676 471 680
rect 475 676 477 680
rect 481 676 483 680
rect 487 676 489 680
rect 493 676 495 680
rect 499 676 509 680
rect 378 674 406 676
rect 382 670 384 674
rect 388 670 390 674
rect 394 670 397 674
rect 401 670 402 674
rect 378 668 406 670
rect 382 664 384 668
rect 388 664 390 668
rect 394 664 397 668
rect 401 664 402 668
rect 378 662 406 664
rect 382 658 384 662
rect 388 658 390 662
rect 394 658 397 662
rect 401 658 402 662
rect 378 656 406 658
rect 382 652 384 656
rect 388 652 390 656
rect 394 652 397 656
rect 401 652 402 656
rect 365 650 369 652
rect 384 650 406 652
rect 388 646 390 650
rect 394 646 397 650
rect 401 646 402 650
rect 413 675 513 676
rect 413 671 414 675
rect 418 671 420 675
rect 424 671 427 675
rect 431 671 433 675
rect 437 671 439 675
rect 443 671 445 675
rect 449 674 513 675
rect 449 671 465 674
rect 413 670 465 671
rect 469 670 471 674
rect 475 670 477 674
rect 481 670 483 674
rect 487 670 489 674
rect 493 670 495 674
rect 499 670 509 674
rect 413 669 513 670
rect 413 665 414 669
rect 418 665 420 669
rect 424 665 427 669
rect 431 665 433 669
rect 437 665 439 669
rect 443 665 445 669
rect 449 668 513 669
rect 449 665 465 668
rect 413 664 465 665
rect 469 664 471 668
rect 475 664 477 668
rect 481 664 483 668
rect 487 664 489 668
rect 493 664 495 668
rect 499 664 509 668
rect 413 663 513 664
rect 413 659 414 663
rect 418 659 420 663
rect 424 659 427 663
rect 431 659 433 663
rect 437 659 439 663
rect 443 659 445 663
rect 449 662 513 663
rect 449 659 465 662
rect 413 658 465 659
rect 469 658 471 662
rect 475 658 477 662
rect 481 658 483 662
rect 487 658 489 662
rect 493 658 495 662
rect 499 658 509 662
rect 413 657 513 658
rect 413 653 414 657
rect 418 653 420 657
rect 424 653 427 657
rect 431 653 433 657
rect 437 653 439 657
rect 443 653 445 657
rect 449 656 513 657
rect 449 653 465 656
rect 413 652 465 653
rect 469 652 471 656
rect 475 652 477 656
rect 481 652 483 656
rect 487 652 489 656
rect 493 652 495 656
rect 499 652 509 656
rect 413 651 513 652
rect 413 647 414 651
rect 418 647 420 651
rect 424 647 427 651
rect 431 647 433 651
rect 437 647 439 651
rect 443 647 445 651
rect 449 650 513 651
rect 449 647 465 650
rect 413 646 465 647
rect 469 646 471 650
rect 475 646 477 650
rect 481 646 483 650
rect 487 646 489 650
rect 493 646 509 650
rect 365 644 369 646
rect 369 640 372 642
rect 365 638 372 640
rect 376 638 412 642
rect 421 638 423 642
rect 427 638 429 642
rect 433 638 435 642
rect 439 638 441 642
rect 450 638 501 642
rect 505 638 509 642
rect 369 636 513 638
rect 369 634 372 636
rect 365 632 372 634
rect 376 632 412 636
rect 421 632 423 636
rect 427 632 429 636
rect 433 632 435 636
rect 439 632 441 636
rect 450 632 501 636
rect 505 632 509 636
rect 369 630 513 632
rect 369 628 372 630
rect 365 626 372 628
rect 376 626 412 630
rect 421 626 423 630
rect 427 626 429 630
rect 433 626 435 630
rect 439 626 441 630
rect 450 626 501 630
rect 505 626 509 630
rect 369 624 513 626
rect 369 622 372 624
rect 365 620 372 622
rect 376 620 412 624
rect 421 620 423 624
rect 427 620 429 624
rect 433 620 435 624
rect 439 620 441 624
rect 450 620 501 624
rect 505 620 509 624
rect 369 618 513 620
rect 369 616 372 618
rect 365 614 372 616
rect 376 614 412 618
rect 421 614 423 618
rect 427 614 429 618
rect 433 614 435 618
rect 439 614 441 618
rect 450 614 501 618
rect 505 614 509 618
rect 369 612 513 614
rect 369 610 372 612
rect 365 608 372 610
rect 376 608 412 612
rect 421 608 423 612
rect 427 608 429 612
rect 433 608 435 612
rect 439 608 441 612
rect 450 608 501 612
rect 505 608 509 612
rect 369 606 513 608
rect 369 604 372 606
rect 365 602 372 604
rect 376 602 412 606
rect 421 602 423 606
rect 427 602 429 606
rect 433 602 435 606
rect 439 602 441 606
rect 450 602 501 606
rect 505 602 509 606
rect 365 596 369 598
rect 365 590 369 592
rect 365 584 369 586
rect 365 578 369 580
rect 365 572 369 574
rect 365 566 369 568
rect 365 560 369 562
rect 365 554 369 556
rect 365 548 369 550
rect 365 542 369 544
rect 365 536 369 538
rect 365 530 369 532
rect 365 524 369 526
rect 365 518 369 520
rect 365 512 369 514
rect 365 506 369 508
rect 365 500 369 502
rect 365 494 369 496
rect 365 488 369 490
rect 365 482 369 484
rect 365 476 369 478
rect 3 472 5 476
rect 9 472 11 476
rect 15 472 17 476
rect 21 472 23 476
rect 27 472 29 476
rect 33 472 35 476
rect 39 472 41 476
rect 45 472 47 476
rect 51 472 53 476
rect 57 472 59 476
rect 63 472 65 476
rect 69 472 71 476
rect 75 472 77 476
rect 81 472 83 476
rect 87 472 89 476
rect 93 472 95 476
rect 99 472 101 476
rect 105 472 107 476
rect 111 472 113 476
rect 117 472 119 476
rect 123 472 125 476
rect 129 472 131 476
rect 135 472 137 476
rect 141 472 143 476
rect 147 472 149 476
rect 153 472 155 476
rect 159 472 161 476
rect 165 472 167 476
rect 171 472 173 476
rect 177 472 179 476
rect 183 472 185 476
rect 189 472 191 476
rect 195 472 197 476
rect 201 472 203 476
rect 207 472 209 476
rect 213 472 215 476
rect 219 472 221 476
rect 225 472 227 476
rect 231 472 233 476
rect 237 472 239 476
rect 243 472 245 476
rect 249 472 251 476
rect 255 472 257 476
rect 261 472 263 476
rect 267 472 269 476
rect 273 472 275 476
rect 279 472 281 476
rect 285 472 287 476
rect 291 472 293 476
rect 297 472 299 476
rect 303 472 305 476
rect 309 472 311 476
rect 315 472 317 476
rect 321 472 323 476
rect 327 472 329 476
rect 333 472 335 476
rect 339 472 341 476
rect 345 472 347 476
rect 351 472 353 476
rect 357 472 359 476
rect 363 472 365 476
rect 365 470 369 472
rect 365 464 369 466
rect 365 458 369 460
rect 365 452 369 454
rect 365 446 369 448
rect 365 440 369 442
rect 365 434 369 436
rect 365 428 369 430
rect 365 422 369 424
rect 365 416 369 418
rect 365 410 369 412
rect 365 404 369 406
rect 365 398 369 400
rect 365 392 369 394
rect 365 386 369 388
rect 365 380 369 382
rect 365 374 369 376
rect 365 368 369 370
rect 365 362 369 364
rect 365 356 369 358
rect 365 350 369 352
rect 365 344 372 346
rect 369 342 372 344
rect 376 342 412 346
rect 421 342 423 346
rect 427 342 429 346
rect 433 342 435 346
rect 439 342 441 346
rect 450 342 501 346
rect 505 342 509 346
rect 369 340 513 342
rect 365 338 372 340
rect 369 336 372 338
rect 376 336 412 340
rect 421 336 423 340
rect 427 336 429 340
rect 433 336 435 340
rect 439 336 441 340
rect 450 336 501 340
rect 505 336 509 340
rect 369 334 513 336
rect 365 332 372 334
rect 369 330 372 332
rect 376 330 412 334
rect 421 330 423 334
rect 427 330 429 334
rect 433 330 435 334
rect 439 330 441 334
rect 450 330 501 334
rect 505 330 509 334
rect 369 328 513 330
rect 365 326 372 328
rect 369 324 372 326
rect 376 324 412 328
rect 421 324 423 328
rect 427 324 429 328
rect 433 324 435 328
rect 439 324 441 328
rect 450 324 501 328
rect 505 324 509 328
rect 369 322 513 324
rect 365 320 372 322
rect 369 318 372 320
rect 376 318 412 322
rect 421 318 423 322
rect 427 318 429 322
rect 433 318 435 322
rect 439 318 441 322
rect 450 318 501 322
rect 505 318 509 322
rect 369 316 513 318
rect 365 314 372 316
rect 369 312 372 314
rect 376 312 412 316
rect 421 312 423 316
rect 427 312 429 316
rect 433 312 435 316
rect 439 312 441 316
rect 450 312 501 316
rect 505 312 509 316
rect 369 310 513 312
rect 365 308 372 310
rect 369 306 372 308
rect 376 306 412 310
rect 421 306 423 310
rect 427 306 429 310
rect 433 306 435 310
rect 439 306 441 310
rect 450 306 501 310
rect 505 306 509 310
rect 365 302 369 304
rect 365 296 369 298
rect 388 298 390 302
rect 394 298 397 302
rect 401 298 402 302
rect 384 296 406 298
rect 365 290 369 292
rect 365 284 369 286
rect 365 278 369 280
rect 365 272 369 274
rect 365 266 369 268
rect 382 292 384 296
rect 388 292 390 296
rect 394 292 397 296
rect 401 292 402 296
rect 378 290 406 292
rect 382 286 384 290
rect 388 286 390 290
rect 394 286 397 290
rect 401 286 402 290
rect 378 284 406 286
rect 382 280 384 284
rect 388 280 390 284
rect 394 280 397 284
rect 401 280 402 284
rect 378 278 406 280
rect 382 274 384 278
rect 388 274 390 278
rect 394 274 397 278
rect 401 274 402 278
rect 378 272 406 274
rect 413 301 465 302
rect 413 297 414 301
rect 418 297 420 301
rect 424 297 427 301
rect 431 297 433 301
rect 437 297 439 301
rect 443 297 445 301
rect 449 298 465 301
rect 469 298 471 302
rect 475 298 477 302
rect 481 298 483 302
rect 487 298 489 302
rect 493 298 509 302
rect 449 297 513 298
rect 413 296 513 297
rect 413 295 465 296
rect 413 291 414 295
rect 418 291 420 295
rect 424 291 427 295
rect 431 291 433 295
rect 437 291 439 295
rect 443 291 445 295
rect 449 292 465 295
rect 469 292 471 296
rect 475 292 477 296
rect 481 292 483 296
rect 487 292 489 296
rect 493 292 495 296
rect 499 292 509 296
rect 449 291 513 292
rect 413 290 513 291
rect 413 289 465 290
rect 413 285 414 289
rect 418 285 420 289
rect 424 285 427 289
rect 431 285 433 289
rect 437 285 439 289
rect 443 285 445 289
rect 449 286 465 289
rect 469 286 471 290
rect 475 286 477 290
rect 481 286 483 290
rect 487 286 489 290
rect 493 286 495 290
rect 499 286 509 290
rect 449 285 513 286
rect 413 284 513 285
rect 413 283 465 284
rect 413 279 414 283
rect 418 279 420 283
rect 424 279 427 283
rect 431 279 433 283
rect 437 279 439 283
rect 443 279 445 283
rect 449 280 465 283
rect 469 280 471 284
rect 475 280 477 284
rect 481 280 483 284
rect 487 280 489 284
rect 493 280 495 284
rect 499 280 509 284
rect 449 279 513 280
rect 413 278 513 279
rect 413 277 465 278
rect 413 273 414 277
rect 418 273 420 277
rect 424 273 427 277
rect 431 273 433 277
rect 437 273 439 277
rect 443 273 445 277
rect 449 274 465 277
rect 469 274 471 278
rect 475 274 477 278
rect 481 274 483 278
rect 487 274 489 278
rect 493 274 495 278
rect 499 274 509 278
rect 449 273 513 274
rect 413 272 513 273
rect 382 268 384 272
rect 388 268 390 272
rect 394 268 397 272
rect 401 268 402 272
rect 469 268 471 272
rect 475 268 477 272
rect 481 268 483 272
rect 487 268 489 272
rect 493 268 495 272
rect 499 268 509 272
rect 378 266 406 268
rect 382 262 384 266
rect 388 262 390 266
rect 394 262 397 266
rect 401 262 402 266
rect 455 264 456 268
rect 460 264 461 268
rect 455 263 461 264
rect 365 260 369 262
rect 365 254 369 256
rect 455 259 456 263
rect 460 259 461 263
rect 465 266 513 268
rect 469 262 471 266
rect 475 262 477 266
rect 481 262 483 266
rect 487 262 489 266
rect 493 262 495 266
rect 499 262 509 266
rect 455 258 461 259
rect 455 254 456 258
rect 460 254 509 258
rect 455 253 509 254
rect 455 249 456 253
rect 460 249 509 253
rect 365 218 369 220
rect 365 212 369 214
rect 455 221 456 225
rect 460 221 509 225
rect 455 220 509 221
rect 455 216 456 220
rect 460 216 509 220
rect 455 215 461 216
rect 365 206 369 208
rect 365 200 369 202
rect 365 194 369 196
rect 365 188 369 190
rect 365 182 369 184
rect 382 208 384 212
rect 388 208 390 212
rect 394 208 397 212
rect 401 208 402 212
rect 378 206 406 208
rect 455 211 456 215
rect 460 211 461 215
rect 455 210 461 211
rect 455 206 456 210
rect 460 206 461 210
rect 469 208 471 212
rect 475 208 477 212
rect 481 208 483 212
rect 487 208 489 212
rect 493 208 495 212
rect 499 208 509 212
rect 465 206 513 208
rect 382 202 384 206
rect 388 202 390 206
rect 394 202 397 206
rect 401 202 402 206
rect 469 202 471 206
rect 475 202 477 206
rect 481 202 483 206
rect 487 202 489 206
rect 493 202 495 206
rect 499 202 509 206
rect 378 200 406 202
rect 382 196 384 200
rect 388 196 390 200
rect 394 196 397 200
rect 401 196 402 200
rect 378 194 406 196
rect 382 190 384 194
rect 388 190 390 194
rect 394 190 397 194
rect 401 190 402 194
rect 378 188 406 190
rect 382 184 384 188
rect 388 184 390 188
rect 394 184 397 188
rect 401 184 402 188
rect 378 182 406 184
rect 382 178 384 182
rect 388 178 390 182
rect 394 178 397 182
rect 401 178 402 182
rect 365 176 369 178
rect 384 176 406 178
rect 388 172 390 176
rect 394 172 397 176
rect 401 172 402 176
rect 413 201 513 202
rect 413 197 414 201
rect 418 197 420 201
rect 424 197 427 201
rect 431 197 433 201
rect 437 197 439 201
rect 443 197 445 201
rect 449 200 513 201
rect 449 197 465 200
rect 413 196 465 197
rect 469 196 471 200
rect 475 196 477 200
rect 481 196 483 200
rect 487 196 489 200
rect 493 196 495 200
rect 499 196 509 200
rect 413 195 513 196
rect 413 191 414 195
rect 418 191 420 195
rect 424 191 427 195
rect 431 191 433 195
rect 437 191 439 195
rect 443 191 445 195
rect 449 194 513 195
rect 449 191 465 194
rect 413 190 465 191
rect 469 190 471 194
rect 475 190 477 194
rect 481 190 483 194
rect 487 190 489 194
rect 493 190 495 194
rect 499 190 509 194
rect 413 189 513 190
rect 413 185 414 189
rect 418 185 420 189
rect 424 185 427 189
rect 431 185 433 189
rect 437 185 439 189
rect 443 185 445 189
rect 449 188 513 189
rect 449 185 465 188
rect 413 184 465 185
rect 469 184 471 188
rect 475 184 477 188
rect 481 184 483 188
rect 487 184 489 188
rect 493 184 495 188
rect 499 184 509 188
rect 413 183 513 184
rect 413 179 414 183
rect 418 179 420 183
rect 424 179 427 183
rect 431 179 433 183
rect 437 179 439 183
rect 443 179 445 183
rect 449 182 513 183
rect 449 179 465 182
rect 413 178 465 179
rect 469 178 471 182
rect 475 178 477 182
rect 481 178 483 182
rect 487 178 489 182
rect 493 178 495 182
rect 499 178 509 182
rect 413 177 513 178
rect 413 173 414 177
rect 418 173 420 177
rect 424 173 427 177
rect 431 173 433 177
rect 437 173 439 177
rect 443 173 445 177
rect 449 176 513 177
rect 449 173 465 176
rect 413 172 465 173
rect 469 172 471 176
rect 475 172 477 176
rect 481 172 483 176
rect 487 172 489 176
rect 493 172 495 176
rect 499 172 509 176
rect 365 170 369 172
rect 369 166 372 168
rect 365 164 372 166
rect 376 164 412 168
rect 421 164 423 168
rect 427 164 429 168
rect 433 164 435 168
rect 439 164 441 168
rect 450 164 451 168
rect 369 162 451 164
rect 369 160 372 162
rect 365 158 372 160
rect 376 158 412 162
rect 421 158 423 162
rect 427 158 429 162
rect 433 158 435 162
rect 439 158 441 162
rect 450 158 451 162
rect 369 156 451 158
rect 369 154 372 156
rect 365 152 372 154
rect 376 152 412 156
rect 421 152 423 156
rect 427 152 429 156
rect 433 152 435 156
rect 439 152 441 156
rect 450 152 451 156
rect 369 150 451 152
rect 369 148 372 150
rect 365 146 372 148
rect 376 146 412 150
rect 421 146 423 150
rect 427 146 429 150
rect 433 146 435 150
rect 439 146 441 150
rect 450 146 451 150
rect 369 144 451 146
rect 369 142 372 144
rect 365 140 372 142
rect 376 140 412 144
rect 421 140 423 144
rect 427 140 429 144
rect 433 140 435 144
rect 439 140 441 144
rect 450 140 451 144
rect 369 138 451 140
rect 369 136 372 138
rect 365 134 372 136
rect 376 134 412 138
rect 421 134 423 138
rect 427 134 429 138
rect 433 134 435 138
rect 439 134 441 138
rect 450 134 451 138
rect 369 132 451 134
rect 369 130 372 132
rect 365 128 372 130
rect 376 128 412 132
rect 421 128 423 132
rect 427 128 429 132
rect 433 128 435 132
rect 439 128 441 132
rect 450 128 451 132
rect 365 122 369 124
rect 365 116 369 118
rect 365 110 369 112
rect 365 104 369 106
rect 365 98 369 100
rect 365 92 369 94
rect 365 86 369 88
rect 365 80 369 82
rect 365 74 369 76
rect 365 68 369 70
rect 365 62 369 64
rect 365 56 369 58
rect 365 50 369 52
rect 365 44 369 46
rect 365 38 369 40
rect 365 32 369 34
rect 365 26 369 28
rect 365 20 369 22
rect 365 14 369 16
rect 365 8 369 10
rect 365 2 369 4
<< m2contact >>
rect 412 4134 421 4138
rect 423 4134 427 4138
rect 429 4134 433 4138
rect 435 4134 439 4138
rect 441 4134 450 4138
rect 412 4128 421 4132
rect 423 4128 427 4132
rect 429 4128 433 4132
rect 435 4128 439 4132
rect 441 4128 450 4132
rect 412 4122 421 4126
rect 423 4122 427 4126
rect 429 4122 433 4126
rect 435 4122 439 4126
rect 441 4122 450 4126
rect 412 4116 421 4120
rect 423 4116 427 4120
rect 429 4116 433 4120
rect 435 4116 439 4120
rect 441 4116 450 4120
rect 412 4110 421 4114
rect 423 4110 427 4114
rect 429 4110 433 4114
rect 435 4110 439 4114
rect 441 4110 450 4114
rect 412 4104 421 4108
rect 423 4104 427 4108
rect 429 4104 433 4108
rect 435 4104 439 4108
rect 441 4104 450 4108
rect 412 4098 421 4102
rect 423 4098 427 4102
rect 429 4098 433 4102
rect 435 4098 439 4102
rect 441 4098 450 4102
rect 390 4090 394 4094
rect 402 4090 406 4094
rect 378 4084 382 4088
rect 390 4084 394 4088
rect 402 4084 406 4088
rect 378 4078 382 4082
rect 390 4078 394 4082
rect 402 4078 406 4082
rect 378 4072 382 4076
rect 390 4072 394 4076
rect 402 4072 406 4076
rect 378 4066 382 4070
rect 390 4066 394 4070
rect 402 4066 406 4070
rect 466 4090 470 4094
rect 477 4090 481 4094
rect 483 4090 487 4094
rect 495 4090 499 4094
rect 509 4090 513 4094
rect 466 4084 470 4088
rect 477 4084 481 4088
rect 483 4084 487 4088
rect 495 4084 499 4088
rect 509 4084 513 4088
rect 466 4078 470 4082
rect 477 4078 481 4082
rect 483 4078 487 4082
rect 495 4078 499 4082
rect 509 4078 513 4082
rect 466 4072 470 4076
rect 477 4072 481 4076
rect 483 4072 487 4076
rect 495 4072 499 4076
rect 509 4072 513 4076
rect 466 4066 470 4070
rect 477 4066 481 4070
rect 483 4066 487 4070
rect 495 4066 499 4070
rect 509 4066 513 4070
rect 378 4060 382 4064
rect 390 4060 394 4064
rect 402 4060 406 4064
rect 466 4060 470 4064
rect 477 4060 481 4064
rect 483 4060 487 4064
rect 495 4060 499 4064
rect 509 4060 513 4064
rect 378 4054 382 4058
rect 390 4054 394 4058
rect 402 4054 406 4058
rect 456 4051 460 4055
rect 466 4054 470 4058
rect 477 4054 481 4058
rect 483 4054 487 4058
rect 495 4054 499 4058
rect 509 4054 513 4058
rect 456 4041 460 4045
rect 509 4041 513 4050
rect 456 4013 460 4017
rect 509 4008 513 4017
rect 378 4000 382 4004
rect 390 4000 394 4004
rect 402 4000 406 4004
rect 456 4003 460 4007
rect 466 4000 470 4004
rect 477 4000 481 4004
rect 483 4000 487 4004
rect 495 4000 499 4004
rect 509 4000 513 4004
rect 378 3994 382 3998
rect 390 3994 394 3998
rect 402 3994 406 3998
rect 466 3994 470 3998
rect 477 3994 481 3998
rect 483 3994 487 3998
rect 495 3994 499 3998
rect 509 3994 513 3998
rect 378 3988 382 3992
rect 390 3988 394 3992
rect 402 3988 406 3992
rect 378 3982 382 3986
rect 390 3982 394 3986
rect 402 3982 406 3986
rect 378 3976 382 3980
rect 390 3976 394 3980
rect 402 3976 406 3980
rect 378 3970 382 3974
rect 390 3970 394 3974
rect 402 3970 406 3974
rect 390 3964 394 3968
rect 402 3964 406 3968
rect 466 3988 470 3992
rect 477 3988 481 3992
rect 483 3988 487 3992
rect 495 3988 499 3992
rect 509 3988 513 3992
rect 466 3982 470 3986
rect 477 3982 481 3986
rect 483 3982 487 3986
rect 495 3982 499 3986
rect 509 3982 513 3986
rect 466 3976 470 3980
rect 477 3976 481 3980
rect 483 3976 487 3980
rect 495 3976 499 3980
rect 509 3976 513 3980
rect 466 3970 470 3974
rect 477 3970 481 3974
rect 483 3970 487 3974
rect 495 3970 499 3974
rect 509 3970 513 3974
rect 466 3964 470 3968
rect 477 3964 481 3968
rect 483 3964 487 3968
rect 509 3964 513 3968
rect 412 3956 421 3960
rect 423 3956 427 3960
rect 429 3956 433 3960
rect 435 3956 439 3960
rect 441 3956 450 3960
rect 509 3956 513 3960
rect 412 3950 421 3954
rect 423 3950 427 3954
rect 429 3950 433 3954
rect 435 3950 439 3954
rect 441 3950 450 3954
rect 509 3950 513 3954
rect 412 3944 421 3948
rect 423 3944 427 3948
rect 429 3944 433 3948
rect 435 3944 439 3948
rect 441 3944 450 3948
rect 509 3944 513 3948
rect 412 3938 421 3942
rect 423 3938 427 3942
rect 429 3938 433 3942
rect 435 3938 439 3942
rect 441 3938 450 3942
rect 509 3938 513 3942
rect 412 3932 421 3936
rect 423 3932 427 3936
rect 429 3932 433 3936
rect 435 3932 439 3936
rect 441 3932 450 3936
rect 509 3932 513 3936
rect 412 3926 421 3930
rect 423 3926 427 3930
rect 429 3926 433 3930
rect 435 3926 439 3930
rect 441 3926 450 3930
rect 509 3926 513 3930
rect 412 3920 421 3924
rect 423 3920 427 3924
rect 429 3920 433 3924
rect 435 3920 439 3924
rect 441 3920 450 3924
rect 509 3920 513 3924
rect 412 3660 421 3664
rect 423 3660 427 3664
rect 429 3660 433 3664
rect 435 3660 439 3664
rect 441 3660 450 3664
rect 509 3660 513 3664
rect 412 3654 421 3658
rect 423 3654 427 3658
rect 429 3654 433 3658
rect 435 3654 439 3658
rect 441 3654 450 3658
rect 509 3654 513 3658
rect 412 3648 421 3652
rect 423 3648 427 3652
rect 429 3648 433 3652
rect 435 3648 439 3652
rect 441 3648 450 3652
rect 509 3648 513 3652
rect 412 3642 421 3646
rect 423 3642 427 3646
rect 429 3642 433 3646
rect 435 3642 439 3646
rect 441 3642 450 3646
rect 509 3642 513 3646
rect 412 3636 421 3640
rect 423 3636 427 3640
rect 429 3636 433 3640
rect 435 3636 439 3640
rect 441 3636 450 3640
rect 509 3636 513 3640
rect 412 3630 421 3634
rect 423 3630 427 3634
rect 429 3630 433 3634
rect 435 3630 439 3634
rect 441 3630 450 3634
rect 509 3630 513 3634
rect 412 3624 421 3628
rect 423 3624 427 3628
rect 429 3624 433 3628
rect 435 3624 439 3628
rect 441 3624 450 3628
rect 509 3624 513 3628
rect 390 3616 394 3620
rect 402 3616 406 3620
rect 378 3610 382 3614
rect 390 3610 394 3614
rect 402 3610 406 3614
rect 378 3604 382 3608
rect 390 3604 394 3608
rect 402 3604 406 3608
rect 378 3598 382 3602
rect 390 3598 394 3602
rect 402 3598 406 3602
rect 378 3592 382 3596
rect 390 3592 394 3596
rect 402 3592 406 3596
rect 465 3616 469 3620
rect 477 3616 481 3620
rect 483 3616 487 3620
rect 509 3616 513 3620
rect 465 3610 469 3614
rect 477 3610 481 3614
rect 483 3610 487 3614
rect 495 3610 499 3614
rect 509 3610 513 3614
rect 465 3604 469 3608
rect 477 3604 481 3608
rect 483 3604 487 3608
rect 495 3604 499 3608
rect 509 3604 513 3608
rect 465 3598 469 3602
rect 477 3598 481 3602
rect 483 3598 487 3602
rect 495 3598 499 3602
rect 509 3598 513 3602
rect 465 3592 469 3596
rect 477 3592 481 3596
rect 483 3592 487 3596
rect 495 3592 499 3596
rect 509 3592 513 3596
rect 378 3586 382 3590
rect 390 3586 394 3590
rect 402 3586 406 3590
rect 465 3586 469 3590
rect 477 3586 481 3590
rect 483 3586 487 3590
rect 495 3586 499 3590
rect 509 3586 513 3590
rect 378 3580 382 3584
rect 390 3580 394 3584
rect 402 3580 406 3584
rect 456 3577 460 3581
rect 465 3580 469 3584
rect 477 3580 481 3584
rect 483 3580 487 3584
rect 495 3580 499 3584
rect 509 3580 513 3584
rect 456 3567 460 3571
rect 509 3567 513 3576
rect 456 3539 460 3543
rect 509 3534 513 3543
rect 378 3526 382 3530
rect 390 3526 394 3530
rect 402 3526 406 3530
rect 456 3529 460 3533
rect 465 3526 469 3530
rect 477 3526 481 3530
rect 483 3526 487 3530
rect 495 3526 499 3530
rect 509 3526 513 3530
rect 378 3520 382 3524
rect 390 3520 394 3524
rect 402 3520 406 3524
rect 465 3520 469 3524
rect 477 3520 481 3524
rect 483 3520 487 3524
rect 495 3520 499 3524
rect 509 3520 513 3524
rect 378 3514 382 3518
rect 390 3514 394 3518
rect 402 3514 406 3518
rect 378 3508 382 3512
rect 390 3508 394 3512
rect 402 3508 406 3512
rect 378 3502 382 3506
rect 390 3502 394 3506
rect 402 3502 406 3506
rect 378 3496 382 3500
rect 390 3496 394 3500
rect 402 3496 406 3500
rect 390 3490 394 3494
rect 402 3490 406 3494
rect 465 3514 469 3518
rect 477 3514 481 3518
rect 483 3514 487 3518
rect 495 3514 499 3518
rect 509 3514 513 3518
rect 465 3508 469 3512
rect 477 3508 481 3512
rect 483 3508 487 3512
rect 495 3508 499 3512
rect 509 3508 513 3512
rect 465 3502 469 3506
rect 477 3502 481 3506
rect 483 3502 487 3506
rect 495 3502 499 3506
rect 509 3502 513 3506
rect 465 3496 469 3500
rect 477 3496 481 3500
rect 483 3496 487 3500
rect 495 3496 499 3500
rect 509 3496 513 3500
rect 465 3490 469 3494
rect 477 3490 481 3494
rect 483 3490 487 3494
rect 509 3490 513 3494
rect 412 3482 421 3486
rect 423 3482 427 3486
rect 429 3482 433 3486
rect 435 3482 439 3486
rect 441 3482 450 3486
rect 509 3482 513 3486
rect 412 3476 421 3480
rect 423 3476 427 3480
rect 429 3476 433 3480
rect 435 3476 439 3480
rect 441 3476 450 3480
rect 509 3476 513 3480
rect 412 3470 421 3474
rect 423 3470 427 3474
rect 429 3470 433 3474
rect 435 3470 439 3474
rect 441 3470 450 3474
rect 509 3470 513 3474
rect 412 3464 421 3468
rect 423 3464 427 3468
rect 429 3464 433 3468
rect 435 3464 439 3468
rect 441 3464 450 3468
rect 509 3464 513 3468
rect 412 3458 421 3462
rect 423 3458 427 3462
rect 429 3458 433 3462
rect 435 3458 439 3462
rect 441 3458 450 3462
rect 509 3458 513 3462
rect 412 3452 421 3456
rect 423 3452 427 3456
rect 429 3452 433 3456
rect 435 3452 439 3456
rect 441 3452 450 3456
rect 509 3452 513 3456
rect 412 3446 421 3450
rect 423 3446 427 3450
rect 429 3446 433 3450
rect 435 3446 439 3450
rect 441 3446 450 3450
rect 509 3446 513 3450
rect 412 3186 421 3190
rect 423 3186 427 3190
rect 429 3186 433 3190
rect 435 3186 439 3190
rect 441 3186 450 3190
rect 509 3186 513 3190
rect 412 3180 421 3184
rect 423 3180 427 3184
rect 429 3180 433 3184
rect 435 3180 439 3184
rect 441 3180 450 3184
rect 509 3180 513 3184
rect 412 3174 421 3178
rect 423 3174 427 3178
rect 429 3174 433 3178
rect 435 3174 439 3178
rect 441 3174 450 3178
rect 509 3174 513 3178
rect 412 3168 421 3172
rect 423 3168 427 3172
rect 429 3168 433 3172
rect 435 3168 439 3172
rect 441 3168 450 3172
rect 509 3168 513 3172
rect 412 3162 421 3166
rect 423 3162 427 3166
rect 429 3162 433 3166
rect 435 3162 439 3166
rect 441 3162 450 3166
rect 509 3162 513 3166
rect 412 3156 421 3160
rect 423 3156 427 3160
rect 429 3156 433 3160
rect 435 3156 439 3160
rect 441 3156 450 3160
rect 509 3156 513 3160
rect 412 3150 421 3154
rect 423 3150 427 3154
rect 429 3150 433 3154
rect 435 3150 439 3154
rect 441 3150 450 3154
rect 509 3150 513 3154
rect 390 3142 394 3146
rect 402 3142 406 3146
rect 378 3136 382 3140
rect 390 3136 394 3140
rect 402 3136 406 3140
rect 378 3130 382 3134
rect 390 3130 394 3134
rect 402 3130 406 3134
rect 378 3124 382 3128
rect 390 3124 394 3128
rect 402 3124 406 3128
rect 378 3118 382 3122
rect 390 3118 394 3122
rect 402 3118 406 3122
rect 465 3142 469 3146
rect 477 3142 481 3146
rect 483 3142 487 3146
rect 509 3142 513 3146
rect 465 3136 469 3140
rect 477 3136 481 3140
rect 483 3136 487 3140
rect 495 3136 499 3140
rect 509 3136 513 3140
rect 465 3130 469 3134
rect 477 3130 481 3134
rect 483 3130 487 3134
rect 495 3130 499 3134
rect 509 3130 513 3134
rect 465 3124 469 3128
rect 477 3124 481 3128
rect 483 3124 487 3128
rect 495 3124 499 3128
rect 509 3124 513 3128
rect 465 3118 469 3122
rect 477 3118 481 3122
rect 483 3118 487 3122
rect 495 3118 499 3122
rect 509 3118 513 3122
rect 378 3112 382 3116
rect 390 3112 394 3116
rect 402 3112 406 3116
rect 465 3112 469 3116
rect 477 3112 481 3116
rect 483 3112 487 3116
rect 495 3112 499 3116
rect 509 3112 513 3116
rect 378 3106 382 3110
rect 390 3106 394 3110
rect 402 3106 406 3110
rect 456 3103 460 3107
rect 465 3106 469 3110
rect 477 3106 481 3110
rect 483 3106 487 3110
rect 495 3106 499 3110
rect 509 3106 513 3110
rect 456 3093 460 3097
rect 509 3093 513 3102
rect 456 3065 460 3069
rect 509 3060 513 3069
rect 378 3052 382 3056
rect 390 3052 394 3056
rect 402 3052 406 3056
rect 456 3055 460 3059
rect 465 3052 469 3056
rect 477 3052 481 3056
rect 483 3052 487 3056
rect 495 3052 499 3056
rect 509 3052 513 3056
rect 378 3046 382 3050
rect 390 3046 394 3050
rect 402 3046 406 3050
rect 465 3046 469 3050
rect 477 3046 481 3050
rect 483 3046 487 3050
rect 495 3046 499 3050
rect 509 3046 513 3050
rect 378 3040 382 3044
rect 390 3040 394 3044
rect 402 3040 406 3044
rect 378 3034 382 3038
rect 390 3034 394 3038
rect 402 3034 406 3038
rect 378 3028 382 3032
rect 390 3028 394 3032
rect 402 3028 406 3032
rect 378 3022 382 3026
rect 390 3022 394 3026
rect 402 3022 406 3026
rect 390 3016 394 3020
rect 402 3016 406 3020
rect 465 3040 469 3044
rect 477 3040 481 3044
rect 483 3040 487 3044
rect 495 3040 499 3044
rect 509 3040 513 3044
rect 465 3034 469 3038
rect 477 3034 481 3038
rect 483 3034 487 3038
rect 495 3034 499 3038
rect 509 3034 513 3038
rect 465 3028 469 3032
rect 477 3028 481 3032
rect 483 3028 487 3032
rect 495 3028 499 3032
rect 509 3028 513 3032
rect 465 3022 469 3026
rect 477 3022 481 3026
rect 483 3022 487 3026
rect 495 3022 499 3026
rect 509 3022 513 3026
rect 465 3016 469 3020
rect 477 3016 481 3020
rect 483 3016 487 3020
rect 509 3016 513 3020
rect 412 3008 421 3012
rect 423 3008 427 3012
rect 429 3008 433 3012
rect 435 3008 439 3012
rect 441 3008 450 3012
rect 509 3008 513 3012
rect 412 3002 421 3006
rect 423 3002 427 3006
rect 429 3002 433 3006
rect 435 3002 439 3006
rect 441 3002 450 3006
rect 509 3002 513 3006
rect 412 2996 421 3000
rect 423 2996 427 3000
rect 429 2996 433 3000
rect 435 2996 439 3000
rect 441 2996 450 3000
rect 509 2996 513 3000
rect 412 2990 421 2994
rect 423 2990 427 2994
rect 429 2990 433 2994
rect 435 2990 439 2994
rect 441 2990 450 2994
rect 509 2990 513 2994
rect 412 2984 421 2988
rect 423 2984 427 2988
rect 429 2984 433 2988
rect 435 2984 439 2988
rect 441 2984 450 2988
rect 509 2984 513 2988
rect 412 2978 421 2982
rect 423 2978 427 2982
rect 429 2978 433 2982
rect 435 2978 439 2982
rect 441 2978 450 2982
rect 509 2978 513 2982
rect 412 2972 421 2976
rect 423 2972 427 2976
rect 429 2972 433 2976
rect 435 2972 439 2976
rect 441 2972 450 2976
rect 509 2972 513 2976
rect 412 2712 421 2716
rect 423 2712 427 2716
rect 429 2712 433 2716
rect 435 2712 439 2716
rect 441 2712 450 2716
rect 509 2712 513 2716
rect 412 2706 421 2710
rect 423 2706 427 2710
rect 429 2706 433 2710
rect 435 2706 439 2710
rect 441 2706 450 2710
rect 509 2706 513 2710
rect 412 2700 421 2704
rect 423 2700 427 2704
rect 429 2700 433 2704
rect 435 2700 439 2704
rect 441 2700 450 2704
rect 509 2700 513 2704
rect 412 2694 421 2698
rect 423 2694 427 2698
rect 429 2694 433 2698
rect 435 2694 439 2698
rect 441 2694 450 2698
rect 509 2694 513 2698
rect 412 2688 421 2692
rect 423 2688 427 2692
rect 429 2688 433 2692
rect 435 2688 439 2692
rect 441 2688 450 2692
rect 509 2688 513 2692
rect 412 2682 421 2686
rect 423 2682 427 2686
rect 429 2682 433 2686
rect 435 2682 439 2686
rect 441 2682 450 2686
rect 509 2682 513 2686
rect 412 2676 421 2680
rect 423 2676 427 2680
rect 429 2676 433 2680
rect 435 2676 439 2680
rect 441 2676 450 2680
rect 509 2676 513 2680
rect 390 2668 394 2672
rect 402 2668 406 2672
rect 378 2662 382 2666
rect 390 2662 394 2666
rect 402 2662 406 2666
rect 378 2656 382 2660
rect 390 2656 394 2660
rect 402 2656 406 2660
rect 378 2650 382 2654
rect 390 2650 394 2654
rect 402 2650 406 2654
rect 378 2644 382 2648
rect 390 2644 394 2648
rect 402 2644 406 2648
rect 465 2668 469 2672
rect 477 2668 481 2672
rect 483 2668 487 2672
rect 509 2668 513 2672
rect 465 2662 469 2666
rect 477 2662 481 2666
rect 483 2662 487 2666
rect 495 2662 499 2666
rect 509 2662 513 2666
rect 465 2656 469 2660
rect 477 2656 481 2660
rect 483 2656 487 2660
rect 495 2656 499 2660
rect 509 2656 513 2660
rect 465 2650 469 2654
rect 477 2650 481 2654
rect 483 2650 487 2654
rect 495 2650 499 2654
rect 509 2650 513 2654
rect 465 2644 469 2648
rect 477 2644 481 2648
rect 483 2644 487 2648
rect 495 2644 499 2648
rect 509 2644 513 2648
rect 378 2638 382 2642
rect 390 2638 394 2642
rect 402 2638 406 2642
rect 465 2638 469 2642
rect 477 2638 481 2642
rect 483 2638 487 2642
rect 495 2638 499 2642
rect 509 2638 513 2642
rect 378 2632 382 2636
rect 390 2632 394 2636
rect 402 2632 406 2636
rect 456 2629 460 2633
rect 465 2632 469 2636
rect 477 2632 481 2636
rect 483 2632 487 2636
rect 495 2632 499 2636
rect 509 2632 513 2636
rect 456 2619 460 2623
rect 509 2619 513 2628
rect 456 2591 460 2595
rect 509 2586 513 2595
rect 378 2578 382 2582
rect 390 2578 394 2582
rect 402 2578 406 2582
rect 456 2581 460 2585
rect 465 2578 469 2582
rect 477 2578 481 2582
rect 483 2578 487 2582
rect 495 2578 499 2582
rect 509 2578 513 2582
rect 378 2572 382 2576
rect 390 2572 394 2576
rect 402 2572 406 2576
rect 465 2572 469 2576
rect 477 2572 481 2576
rect 483 2572 487 2576
rect 495 2572 499 2576
rect 509 2572 513 2576
rect 378 2566 382 2570
rect 390 2566 394 2570
rect 402 2566 406 2570
rect 378 2560 382 2564
rect 390 2560 394 2564
rect 402 2560 406 2564
rect 378 2554 382 2558
rect 390 2554 394 2558
rect 402 2554 406 2558
rect 378 2548 382 2552
rect 390 2548 394 2552
rect 402 2548 406 2552
rect 390 2542 394 2546
rect 402 2542 406 2546
rect 465 2566 469 2570
rect 477 2566 481 2570
rect 483 2566 487 2570
rect 495 2566 499 2570
rect 509 2566 513 2570
rect 465 2560 469 2564
rect 477 2560 481 2564
rect 483 2560 487 2564
rect 495 2560 499 2564
rect 509 2560 513 2564
rect 465 2554 469 2558
rect 477 2554 481 2558
rect 483 2554 487 2558
rect 495 2554 499 2558
rect 509 2554 513 2558
rect 465 2548 469 2552
rect 477 2548 481 2552
rect 483 2548 487 2552
rect 495 2548 499 2552
rect 509 2548 513 2552
rect 465 2542 469 2546
rect 477 2542 481 2546
rect 483 2542 487 2546
rect 509 2542 513 2546
rect 412 2534 421 2538
rect 423 2534 427 2538
rect 429 2534 433 2538
rect 435 2534 439 2538
rect 441 2534 450 2538
rect 509 2534 513 2538
rect 412 2528 421 2532
rect 423 2528 427 2532
rect 429 2528 433 2532
rect 435 2528 439 2532
rect 441 2528 450 2532
rect 509 2528 513 2532
rect 412 2522 421 2526
rect 423 2522 427 2526
rect 429 2522 433 2526
rect 435 2522 439 2526
rect 441 2522 450 2526
rect 509 2522 513 2526
rect 412 2516 421 2520
rect 423 2516 427 2520
rect 429 2516 433 2520
rect 435 2516 439 2520
rect 441 2516 450 2520
rect 509 2516 513 2520
rect 412 2510 421 2514
rect 423 2510 427 2514
rect 429 2510 433 2514
rect 435 2510 439 2514
rect 441 2510 450 2514
rect 509 2510 513 2514
rect 412 2504 421 2508
rect 423 2504 427 2508
rect 429 2504 433 2508
rect 435 2504 439 2508
rect 441 2504 450 2508
rect 509 2504 513 2508
rect 412 2498 421 2502
rect 423 2498 427 2502
rect 429 2498 433 2502
rect 435 2498 439 2502
rect 441 2498 450 2502
rect 509 2498 513 2502
rect 412 2238 421 2242
rect 423 2238 427 2242
rect 429 2238 433 2242
rect 435 2238 439 2242
rect 441 2238 450 2242
rect 509 2238 513 2242
rect 412 2232 421 2236
rect 423 2232 427 2236
rect 429 2232 433 2236
rect 435 2232 439 2236
rect 441 2232 450 2236
rect 509 2232 513 2236
rect 412 2226 421 2230
rect 423 2226 427 2230
rect 429 2226 433 2230
rect 435 2226 439 2230
rect 441 2226 450 2230
rect 509 2226 513 2230
rect 412 2220 421 2224
rect 423 2220 427 2224
rect 429 2220 433 2224
rect 435 2220 439 2224
rect 441 2220 450 2224
rect 509 2220 513 2224
rect 412 2214 421 2218
rect 423 2214 427 2218
rect 429 2214 433 2218
rect 435 2214 439 2218
rect 441 2214 450 2218
rect 509 2214 513 2218
rect 412 2208 421 2212
rect 423 2208 427 2212
rect 429 2208 433 2212
rect 435 2208 439 2212
rect 441 2208 450 2212
rect 509 2208 513 2212
rect 412 2202 421 2206
rect 423 2202 427 2206
rect 429 2202 433 2206
rect 435 2202 439 2206
rect 441 2202 450 2206
rect 509 2202 513 2206
rect 390 2194 394 2198
rect 402 2194 406 2198
rect 378 2188 382 2192
rect 390 2188 394 2192
rect 402 2188 406 2192
rect 378 2182 382 2186
rect 390 2182 394 2186
rect 402 2182 406 2186
rect 378 2176 382 2180
rect 390 2176 394 2180
rect 402 2176 406 2180
rect 378 2170 382 2174
rect 390 2170 394 2174
rect 402 2170 406 2174
rect 465 2194 469 2198
rect 477 2194 481 2198
rect 483 2194 487 2198
rect 509 2194 513 2198
rect 465 2188 469 2192
rect 477 2188 481 2192
rect 483 2188 487 2192
rect 495 2188 499 2192
rect 509 2188 513 2192
rect 465 2182 469 2186
rect 477 2182 481 2186
rect 483 2182 487 2186
rect 495 2182 499 2186
rect 509 2182 513 2186
rect 465 2176 469 2180
rect 477 2176 481 2180
rect 483 2176 487 2180
rect 495 2176 499 2180
rect 509 2176 513 2180
rect 465 2170 469 2174
rect 477 2170 481 2174
rect 483 2170 487 2174
rect 495 2170 499 2174
rect 509 2170 513 2174
rect 378 2164 382 2168
rect 390 2164 394 2168
rect 402 2164 406 2168
rect 465 2164 469 2168
rect 477 2164 481 2168
rect 483 2164 487 2168
rect 495 2164 499 2168
rect 509 2164 513 2168
rect 378 2158 382 2162
rect 390 2158 394 2162
rect 402 2158 406 2162
rect 456 2155 460 2159
rect 465 2158 469 2162
rect 477 2158 481 2162
rect 483 2158 487 2162
rect 495 2158 499 2162
rect 509 2158 513 2162
rect 456 2145 460 2149
rect 509 2145 513 2154
rect 456 2117 460 2121
rect 509 2112 513 2121
rect 378 2104 382 2108
rect 390 2104 394 2108
rect 402 2104 406 2108
rect 456 2107 460 2111
rect 465 2104 469 2108
rect 477 2104 481 2108
rect 483 2104 487 2108
rect 495 2104 499 2108
rect 509 2104 513 2108
rect 378 2098 382 2102
rect 390 2098 394 2102
rect 402 2098 406 2102
rect 465 2098 469 2102
rect 477 2098 481 2102
rect 483 2098 487 2102
rect 495 2098 499 2102
rect 509 2098 513 2102
rect 378 2092 382 2096
rect 390 2092 394 2096
rect 402 2092 406 2096
rect 378 2086 382 2090
rect 390 2086 394 2090
rect 402 2086 406 2090
rect 378 2080 382 2084
rect 390 2080 394 2084
rect 402 2080 406 2084
rect 378 2074 382 2078
rect 390 2074 394 2078
rect 402 2074 406 2078
rect 390 2068 394 2072
rect 402 2068 406 2072
rect 465 2092 469 2096
rect 477 2092 481 2096
rect 483 2092 487 2096
rect 495 2092 499 2096
rect 509 2092 513 2096
rect 465 2086 469 2090
rect 477 2086 481 2090
rect 483 2086 487 2090
rect 495 2086 499 2090
rect 509 2086 513 2090
rect 465 2080 469 2084
rect 477 2080 481 2084
rect 483 2080 487 2084
rect 495 2080 499 2084
rect 509 2080 513 2084
rect 465 2074 469 2078
rect 477 2074 481 2078
rect 483 2074 487 2078
rect 495 2074 499 2078
rect 509 2074 513 2078
rect 465 2068 469 2072
rect 477 2068 481 2072
rect 483 2068 487 2072
rect 509 2068 513 2072
rect 412 2060 421 2064
rect 423 2060 427 2064
rect 429 2060 433 2064
rect 435 2060 439 2064
rect 441 2060 450 2064
rect 509 2060 513 2064
rect 412 2054 421 2058
rect 423 2054 427 2058
rect 429 2054 433 2058
rect 435 2054 439 2058
rect 441 2054 450 2058
rect 509 2054 513 2058
rect 412 2048 421 2052
rect 423 2048 427 2052
rect 429 2048 433 2052
rect 435 2048 439 2052
rect 441 2048 450 2052
rect 509 2048 513 2052
rect 412 2042 421 2046
rect 423 2042 427 2046
rect 429 2042 433 2046
rect 435 2042 439 2046
rect 441 2042 450 2046
rect 509 2042 513 2046
rect 412 2036 421 2040
rect 423 2036 427 2040
rect 429 2036 433 2040
rect 435 2036 439 2040
rect 441 2036 450 2040
rect 509 2036 513 2040
rect 412 2030 421 2034
rect 423 2030 427 2034
rect 429 2030 433 2034
rect 435 2030 439 2034
rect 441 2030 450 2034
rect 509 2030 513 2034
rect 412 2024 421 2028
rect 423 2024 427 2028
rect 429 2024 433 2028
rect 435 2024 439 2028
rect 441 2024 450 2028
rect 509 2024 513 2028
rect 412 1764 421 1768
rect 423 1764 427 1768
rect 429 1764 433 1768
rect 435 1764 439 1768
rect 441 1764 450 1768
rect 509 1764 513 1768
rect 412 1758 421 1762
rect 423 1758 427 1762
rect 429 1758 433 1762
rect 435 1758 439 1762
rect 441 1758 450 1762
rect 509 1758 513 1762
rect 412 1752 421 1756
rect 423 1752 427 1756
rect 429 1752 433 1756
rect 435 1752 439 1756
rect 441 1752 450 1756
rect 509 1752 513 1756
rect 412 1746 421 1750
rect 423 1746 427 1750
rect 429 1746 433 1750
rect 435 1746 439 1750
rect 441 1746 450 1750
rect 509 1746 513 1750
rect 412 1740 421 1744
rect 423 1740 427 1744
rect 429 1740 433 1744
rect 435 1740 439 1744
rect 441 1740 450 1744
rect 509 1740 513 1744
rect 412 1734 421 1738
rect 423 1734 427 1738
rect 429 1734 433 1738
rect 435 1734 439 1738
rect 441 1734 450 1738
rect 509 1734 513 1738
rect 412 1728 421 1732
rect 423 1728 427 1732
rect 429 1728 433 1732
rect 435 1728 439 1732
rect 441 1728 450 1732
rect 509 1728 513 1732
rect 390 1720 394 1724
rect 402 1720 406 1724
rect 378 1714 382 1718
rect 390 1714 394 1718
rect 402 1714 406 1718
rect 378 1708 382 1712
rect 390 1708 394 1712
rect 402 1708 406 1712
rect 378 1702 382 1706
rect 390 1702 394 1706
rect 402 1702 406 1706
rect 378 1696 382 1700
rect 390 1696 394 1700
rect 402 1696 406 1700
rect 465 1720 469 1724
rect 477 1720 481 1724
rect 483 1720 487 1724
rect 509 1720 513 1724
rect 465 1714 469 1718
rect 477 1714 481 1718
rect 483 1714 487 1718
rect 495 1714 499 1718
rect 509 1714 513 1718
rect 465 1708 469 1712
rect 477 1708 481 1712
rect 483 1708 487 1712
rect 495 1708 499 1712
rect 509 1708 513 1712
rect 465 1702 469 1706
rect 477 1702 481 1706
rect 483 1702 487 1706
rect 495 1702 499 1706
rect 509 1702 513 1706
rect 465 1696 469 1700
rect 477 1696 481 1700
rect 483 1696 487 1700
rect 495 1696 499 1700
rect 509 1696 513 1700
rect 378 1690 382 1694
rect 390 1690 394 1694
rect 402 1690 406 1694
rect 465 1690 469 1694
rect 477 1690 481 1694
rect 483 1690 487 1694
rect 495 1690 499 1694
rect 509 1690 513 1694
rect 378 1684 382 1688
rect 390 1684 394 1688
rect 402 1684 406 1688
rect 456 1681 460 1685
rect 465 1684 469 1688
rect 477 1684 481 1688
rect 483 1684 487 1688
rect 495 1684 499 1688
rect 509 1684 513 1688
rect 456 1671 460 1675
rect 509 1671 513 1680
rect 456 1643 460 1647
rect 509 1638 513 1647
rect 378 1630 382 1634
rect 390 1630 394 1634
rect 402 1630 406 1634
rect 456 1633 460 1637
rect 465 1630 469 1634
rect 477 1630 481 1634
rect 483 1630 487 1634
rect 495 1630 499 1634
rect 509 1630 513 1634
rect 378 1624 382 1628
rect 390 1624 394 1628
rect 402 1624 406 1628
rect 465 1624 469 1628
rect 477 1624 481 1628
rect 483 1624 487 1628
rect 495 1624 499 1628
rect 509 1624 513 1628
rect 378 1618 382 1622
rect 390 1618 394 1622
rect 402 1618 406 1622
rect 378 1612 382 1616
rect 390 1612 394 1616
rect 402 1612 406 1616
rect 378 1606 382 1610
rect 390 1606 394 1610
rect 402 1606 406 1610
rect 378 1600 382 1604
rect 390 1600 394 1604
rect 402 1600 406 1604
rect 390 1594 394 1598
rect 402 1594 406 1598
rect 465 1618 469 1622
rect 477 1618 481 1622
rect 483 1618 487 1622
rect 495 1618 499 1622
rect 509 1618 513 1622
rect 465 1612 469 1616
rect 477 1612 481 1616
rect 483 1612 487 1616
rect 495 1612 499 1616
rect 509 1612 513 1616
rect 465 1606 469 1610
rect 477 1606 481 1610
rect 483 1606 487 1610
rect 495 1606 499 1610
rect 509 1606 513 1610
rect 465 1600 469 1604
rect 477 1600 481 1604
rect 483 1600 487 1604
rect 495 1600 499 1604
rect 509 1600 513 1604
rect 465 1594 469 1598
rect 477 1594 481 1598
rect 483 1594 487 1598
rect 509 1594 513 1598
rect 412 1586 421 1590
rect 423 1586 427 1590
rect 429 1586 433 1590
rect 435 1586 439 1590
rect 441 1586 450 1590
rect 509 1586 513 1590
rect 412 1580 421 1584
rect 423 1580 427 1584
rect 429 1580 433 1584
rect 435 1580 439 1584
rect 441 1580 450 1584
rect 509 1580 513 1584
rect 412 1574 421 1578
rect 423 1574 427 1578
rect 429 1574 433 1578
rect 435 1574 439 1578
rect 441 1574 450 1578
rect 509 1574 513 1578
rect 412 1568 421 1572
rect 423 1568 427 1572
rect 429 1568 433 1572
rect 435 1568 439 1572
rect 441 1568 450 1572
rect 509 1568 513 1572
rect 412 1562 421 1566
rect 423 1562 427 1566
rect 429 1562 433 1566
rect 435 1562 439 1566
rect 441 1562 450 1566
rect 509 1562 513 1566
rect 412 1556 421 1560
rect 423 1556 427 1560
rect 429 1556 433 1560
rect 435 1556 439 1560
rect 441 1556 450 1560
rect 509 1556 513 1560
rect 412 1550 421 1554
rect 423 1550 427 1554
rect 429 1550 433 1554
rect 435 1550 439 1554
rect 441 1550 450 1554
rect 509 1550 513 1554
rect 412 1290 421 1294
rect 423 1290 427 1294
rect 429 1290 433 1294
rect 435 1290 439 1294
rect 441 1290 450 1294
rect 509 1290 513 1294
rect 412 1284 421 1288
rect 423 1284 427 1288
rect 429 1284 433 1288
rect 435 1284 439 1288
rect 441 1284 450 1288
rect 509 1284 513 1288
rect 412 1278 421 1282
rect 423 1278 427 1282
rect 429 1278 433 1282
rect 435 1278 439 1282
rect 441 1278 450 1282
rect 509 1278 513 1282
rect 412 1272 421 1276
rect 423 1272 427 1276
rect 429 1272 433 1276
rect 435 1272 439 1276
rect 441 1272 450 1276
rect 509 1272 513 1276
rect 412 1266 421 1270
rect 423 1266 427 1270
rect 429 1266 433 1270
rect 435 1266 439 1270
rect 441 1266 450 1270
rect 509 1266 513 1270
rect 412 1260 421 1264
rect 423 1260 427 1264
rect 429 1260 433 1264
rect 435 1260 439 1264
rect 441 1260 450 1264
rect 509 1260 513 1264
rect 412 1254 421 1258
rect 423 1254 427 1258
rect 429 1254 433 1258
rect 435 1254 439 1258
rect 441 1254 450 1258
rect 509 1254 513 1258
rect 390 1246 394 1250
rect 402 1246 406 1250
rect 378 1240 382 1244
rect 390 1240 394 1244
rect 402 1240 406 1244
rect 378 1234 382 1238
rect 390 1234 394 1238
rect 402 1234 406 1238
rect 378 1228 382 1232
rect 390 1228 394 1232
rect 402 1228 406 1232
rect 378 1222 382 1226
rect 390 1222 394 1226
rect 402 1222 406 1226
rect 465 1246 469 1250
rect 477 1246 481 1250
rect 483 1246 487 1250
rect 509 1246 513 1250
rect 465 1240 469 1244
rect 477 1240 481 1244
rect 483 1240 487 1244
rect 495 1240 499 1244
rect 509 1240 513 1244
rect 465 1234 469 1238
rect 477 1234 481 1238
rect 483 1234 487 1238
rect 495 1234 499 1238
rect 509 1234 513 1238
rect 465 1228 469 1232
rect 477 1228 481 1232
rect 483 1228 487 1232
rect 495 1228 499 1232
rect 509 1228 513 1232
rect 465 1222 469 1226
rect 477 1222 481 1226
rect 483 1222 487 1226
rect 495 1222 499 1226
rect 509 1222 513 1226
rect 378 1216 382 1220
rect 390 1216 394 1220
rect 402 1216 406 1220
rect 465 1216 469 1220
rect 477 1216 481 1220
rect 483 1216 487 1220
rect 495 1216 499 1220
rect 509 1216 513 1220
rect 378 1210 382 1214
rect 390 1210 394 1214
rect 402 1210 406 1214
rect 456 1207 460 1211
rect 465 1210 469 1214
rect 477 1210 481 1214
rect 483 1210 487 1214
rect 495 1210 499 1214
rect 509 1210 513 1214
rect 456 1197 460 1201
rect 509 1197 513 1206
rect 456 1169 460 1173
rect 509 1164 513 1173
rect 378 1156 382 1160
rect 390 1156 394 1160
rect 402 1156 406 1160
rect 456 1159 460 1163
rect 465 1156 469 1160
rect 477 1156 481 1160
rect 483 1156 487 1160
rect 495 1156 499 1160
rect 509 1156 513 1160
rect 378 1150 382 1154
rect 390 1150 394 1154
rect 402 1150 406 1154
rect 465 1150 469 1154
rect 477 1150 481 1154
rect 483 1150 487 1154
rect 495 1150 499 1154
rect 509 1150 513 1154
rect 378 1144 382 1148
rect 390 1144 394 1148
rect 402 1144 406 1148
rect 378 1138 382 1142
rect 390 1138 394 1142
rect 402 1138 406 1142
rect 378 1132 382 1136
rect 390 1132 394 1136
rect 402 1132 406 1136
rect 378 1126 382 1130
rect 390 1126 394 1130
rect 402 1126 406 1130
rect 390 1120 394 1124
rect 402 1120 406 1124
rect 465 1144 469 1148
rect 477 1144 481 1148
rect 483 1144 487 1148
rect 495 1144 499 1148
rect 509 1144 513 1148
rect 465 1138 469 1142
rect 477 1138 481 1142
rect 483 1138 487 1142
rect 495 1138 499 1142
rect 509 1138 513 1142
rect 465 1132 469 1136
rect 477 1132 481 1136
rect 483 1132 487 1136
rect 495 1132 499 1136
rect 509 1132 513 1136
rect 465 1126 469 1130
rect 477 1126 481 1130
rect 483 1126 487 1130
rect 495 1126 499 1130
rect 509 1126 513 1130
rect 465 1120 469 1124
rect 477 1120 481 1124
rect 483 1120 487 1124
rect 509 1120 513 1124
rect 412 1112 421 1116
rect 423 1112 427 1116
rect 429 1112 433 1116
rect 435 1112 439 1116
rect 441 1112 450 1116
rect 509 1112 513 1116
rect 412 1106 421 1110
rect 423 1106 427 1110
rect 429 1106 433 1110
rect 435 1106 439 1110
rect 441 1106 450 1110
rect 509 1106 513 1110
rect 412 1100 421 1104
rect 423 1100 427 1104
rect 429 1100 433 1104
rect 435 1100 439 1104
rect 441 1100 450 1104
rect 509 1100 513 1104
rect 412 1094 421 1098
rect 423 1094 427 1098
rect 429 1094 433 1098
rect 435 1094 439 1098
rect 441 1094 450 1098
rect 509 1094 513 1098
rect 412 1088 421 1092
rect 423 1088 427 1092
rect 429 1088 433 1092
rect 435 1088 439 1092
rect 441 1088 450 1092
rect 509 1088 513 1092
rect 412 1082 421 1086
rect 423 1082 427 1086
rect 429 1082 433 1086
rect 435 1082 439 1086
rect 441 1082 450 1086
rect 509 1082 513 1086
rect 412 1076 421 1080
rect 423 1076 427 1080
rect 429 1076 433 1080
rect 435 1076 439 1080
rect 441 1076 450 1080
rect 509 1076 513 1080
rect 412 816 421 820
rect 423 816 427 820
rect 429 816 433 820
rect 435 816 439 820
rect 441 816 450 820
rect 509 816 513 820
rect 412 810 421 814
rect 423 810 427 814
rect 429 810 433 814
rect 435 810 439 814
rect 441 810 450 814
rect 509 810 513 814
rect 412 804 421 808
rect 423 804 427 808
rect 429 804 433 808
rect 435 804 439 808
rect 441 804 450 808
rect 509 804 513 808
rect 412 798 421 802
rect 423 798 427 802
rect 429 798 433 802
rect 435 798 439 802
rect 441 798 450 802
rect 509 798 513 802
rect 412 792 421 796
rect 423 792 427 796
rect 429 792 433 796
rect 435 792 439 796
rect 441 792 450 796
rect 509 792 513 796
rect 412 786 421 790
rect 423 786 427 790
rect 429 786 433 790
rect 435 786 439 790
rect 441 786 450 790
rect 509 786 513 790
rect 412 780 421 784
rect 423 780 427 784
rect 429 780 433 784
rect 435 780 439 784
rect 441 780 450 784
rect 509 780 513 784
rect 390 772 394 776
rect 402 772 406 776
rect 378 766 382 770
rect 390 766 394 770
rect 402 766 406 770
rect 378 760 382 764
rect 390 760 394 764
rect 402 760 406 764
rect 378 754 382 758
rect 390 754 394 758
rect 402 754 406 758
rect 378 748 382 752
rect 390 748 394 752
rect 402 748 406 752
rect 465 772 469 776
rect 477 772 481 776
rect 483 772 487 776
rect 509 772 513 776
rect 465 766 469 770
rect 477 766 481 770
rect 483 766 487 770
rect 495 766 499 770
rect 509 766 513 770
rect 465 760 469 764
rect 477 760 481 764
rect 483 760 487 764
rect 495 760 499 764
rect 509 760 513 764
rect 465 754 469 758
rect 477 754 481 758
rect 483 754 487 758
rect 495 754 499 758
rect 509 754 513 758
rect 465 748 469 752
rect 477 748 481 752
rect 483 748 487 752
rect 495 748 499 752
rect 509 748 513 752
rect 378 742 382 746
rect 390 742 394 746
rect 402 742 406 746
rect 465 742 469 746
rect 477 742 481 746
rect 483 742 487 746
rect 495 742 499 746
rect 509 742 513 746
rect 378 736 382 740
rect 390 736 394 740
rect 402 736 406 740
rect 456 733 460 737
rect 465 736 469 740
rect 477 736 481 740
rect 483 736 487 740
rect 495 736 499 740
rect 509 736 513 740
rect 456 723 460 727
rect 509 723 513 732
rect 456 695 460 699
rect 509 690 513 699
rect 378 682 382 686
rect 390 682 394 686
rect 402 682 406 686
rect 456 685 460 689
rect 465 682 469 686
rect 477 682 481 686
rect 483 682 487 686
rect 495 682 499 686
rect 509 682 513 686
rect 378 676 382 680
rect 390 676 394 680
rect 402 676 406 680
rect 465 676 469 680
rect 477 676 481 680
rect 483 676 487 680
rect 495 676 499 680
rect 509 676 513 680
rect 378 670 382 674
rect 390 670 394 674
rect 402 670 406 674
rect 378 664 382 668
rect 390 664 394 668
rect 402 664 406 668
rect 378 658 382 662
rect 390 658 394 662
rect 402 658 406 662
rect 378 652 382 656
rect 390 652 394 656
rect 402 652 406 656
rect 390 646 394 650
rect 402 646 406 650
rect 465 670 469 674
rect 477 670 481 674
rect 483 670 487 674
rect 495 670 499 674
rect 509 670 513 674
rect 465 664 469 668
rect 477 664 481 668
rect 483 664 487 668
rect 495 664 499 668
rect 509 664 513 668
rect 465 658 469 662
rect 477 658 481 662
rect 483 658 487 662
rect 495 658 499 662
rect 509 658 513 662
rect 465 652 469 656
rect 477 652 481 656
rect 483 652 487 656
rect 495 652 499 656
rect 509 652 513 656
rect 465 646 469 650
rect 477 646 481 650
rect 483 646 487 650
rect 509 646 513 650
rect 412 638 421 642
rect 423 638 427 642
rect 429 638 433 642
rect 435 638 439 642
rect 441 638 450 642
rect 509 638 513 642
rect 412 632 421 636
rect 423 632 427 636
rect 429 632 433 636
rect 435 632 439 636
rect 441 632 450 636
rect 509 632 513 636
rect 412 626 421 630
rect 423 626 427 630
rect 429 626 433 630
rect 435 626 439 630
rect 441 626 450 630
rect 509 626 513 630
rect 412 620 421 624
rect 423 620 427 624
rect 429 620 433 624
rect 435 620 439 624
rect 441 620 450 624
rect 509 620 513 624
rect 412 614 421 618
rect 423 614 427 618
rect 429 614 433 618
rect 435 614 439 618
rect 441 614 450 618
rect 509 614 513 618
rect 412 608 421 612
rect 423 608 427 612
rect 429 608 433 612
rect 435 608 439 612
rect 441 608 450 612
rect 509 608 513 612
rect 412 602 421 606
rect 423 602 427 606
rect 429 602 433 606
rect 435 602 439 606
rect 441 602 450 606
rect 509 602 513 606
rect 412 342 421 346
rect 423 342 427 346
rect 429 342 433 346
rect 435 342 439 346
rect 441 342 450 346
rect 509 342 513 346
rect 412 336 421 340
rect 423 336 427 340
rect 429 336 433 340
rect 435 336 439 340
rect 441 336 450 340
rect 509 336 513 340
rect 412 330 421 334
rect 423 330 427 334
rect 429 330 433 334
rect 435 330 439 334
rect 441 330 450 334
rect 509 330 513 334
rect 412 324 421 328
rect 423 324 427 328
rect 429 324 433 328
rect 435 324 439 328
rect 441 324 450 328
rect 509 324 513 328
rect 412 318 421 322
rect 423 318 427 322
rect 429 318 433 322
rect 435 318 439 322
rect 441 318 450 322
rect 509 318 513 322
rect 412 312 421 316
rect 423 312 427 316
rect 429 312 433 316
rect 435 312 439 316
rect 441 312 450 316
rect 509 312 513 316
rect 412 306 421 310
rect 423 306 427 310
rect 429 306 433 310
rect 435 306 439 310
rect 441 306 450 310
rect 509 306 513 310
rect 390 298 394 302
rect 402 298 406 302
rect 378 292 382 296
rect 390 292 394 296
rect 402 292 406 296
rect 378 286 382 290
rect 390 286 394 290
rect 402 286 406 290
rect 378 280 382 284
rect 390 280 394 284
rect 402 280 406 284
rect 378 274 382 278
rect 390 274 394 278
rect 402 274 406 278
rect 465 298 469 302
rect 477 298 481 302
rect 483 298 487 302
rect 509 298 513 302
rect 465 292 469 296
rect 477 292 481 296
rect 483 292 487 296
rect 495 292 499 296
rect 509 292 513 296
rect 465 286 469 290
rect 477 286 481 290
rect 483 286 487 290
rect 495 286 499 290
rect 509 286 513 290
rect 465 280 469 284
rect 477 280 481 284
rect 483 280 487 284
rect 495 280 499 284
rect 509 280 513 284
rect 465 274 469 278
rect 477 274 481 278
rect 483 274 487 278
rect 495 274 499 278
rect 509 274 513 278
rect 378 268 382 272
rect 390 268 394 272
rect 402 268 406 272
rect 465 268 469 272
rect 477 268 481 272
rect 483 268 487 272
rect 495 268 499 272
rect 509 268 513 272
rect 378 262 382 266
rect 390 262 394 266
rect 402 262 406 266
rect 456 259 460 263
rect 465 262 469 266
rect 477 262 481 266
rect 483 262 487 266
rect 495 262 499 266
rect 509 262 513 266
rect 456 249 460 253
rect 509 249 513 258
rect 456 221 460 225
rect 509 216 513 225
rect 378 208 382 212
rect 390 208 394 212
rect 402 208 406 212
rect 456 211 460 215
rect 465 208 469 212
rect 477 208 481 212
rect 483 208 487 212
rect 495 208 499 212
rect 509 208 513 212
rect 378 202 382 206
rect 390 202 394 206
rect 402 202 406 206
rect 465 202 469 206
rect 477 202 481 206
rect 483 202 487 206
rect 495 202 499 206
rect 509 202 513 206
rect 378 196 382 200
rect 390 196 394 200
rect 402 196 406 200
rect 378 190 382 194
rect 390 190 394 194
rect 402 190 406 194
rect 378 184 382 188
rect 390 184 394 188
rect 402 184 406 188
rect 378 178 382 182
rect 390 178 394 182
rect 402 178 406 182
rect 390 172 394 176
rect 402 172 406 176
rect 465 196 469 200
rect 477 196 481 200
rect 483 196 487 200
rect 495 196 499 200
rect 509 196 513 200
rect 465 190 469 194
rect 477 190 481 194
rect 483 190 487 194
rect 495 190 499 194
rect 509 190 513 194
rect 465 184 469 188
rect 477 184 481 188
rect 483 184 487 188
rect 495 184 499 188
rect 509 184 513 188
rect 465 178 469 182
rect 477 178 481 182
rect 483 178 487 182
rect 495 178 499 182
rect 509 178 513 182
rect 465 172 469 176
rect 477 172 481 176
rect 483 172 487 176
rect 495 172 499 176
rect 509 172 513 176
rect 412 164 421 168
rect 423 164 427 168
rect 429 164 433 168
rect 435 164 439 168
rect 441 164 450 168
rect 412 158 421 162
rect 423 158 427 162
rect 429 158 433 162
rect 435 158 439 162
rect 441 158 450 162
rect 412 152 421 156
rect 423 152 427 156
rect 429 152 433 156
rect 435 152 439 156
rect 441 152 450 156
rect 412 146 421 150
rect 423 146 427 150
rect 429 146 433 150
rect 435 146 439 150
rect 441 146 450 150
rect 412 140 421 144
rect 423 140 427 144
rect 429 140 433 144
rect 435 140 439 144
rect 441 140 450 144
rect 412 134 421 138
rect 423 134 427 138
rect 429 134 433 138
rect 435 134 439 138
rect 441 134 450 138
rect 412 128 421 132
rect 423 128 427 132
rect 429 128 433 132
rect 435 128 439 132
rect 441 128 450 132
<< metal2 >>
rect 367 4094 407 4226
rect 367 4090 390 4094
rect 394 4090 402 4094
rect 406 4090 407 4094
rect 367 4088 407 4090
rect 367 4084 378 4088
rect 382 4084 390 4088
rect 394 4084 402 4088
rect 406 4084 407 4088
rect 367 4082 407 4084
rect 367 4078 378 4082
rect 382 4078 390 4082
rect 394 4078 402 4082
rect 406 4078 407 4082
rect 367 4076 407 4078
rect 367 4072 378 4076
rect 382 4072 390 4076
rect 394 4072 402 4076
rect 406 4072 407 4076
rect 367 4070 407 4072
rect 367 4066 378 4070
rect 382 4066 390 4070
rect 394 4066 402 4070
rect 406 4066 407 4070
rect 367 4064 407 4066
rect 367 4060 378 4064
rect 382 4060 390 4064
rect 394 4060 402 4064
rect 406 4060 407 4064
rect 367 4058 407 4060
rect 367 4054 378 4058
rect 382 4054 390 4058
rect 394 4054 402 4058
rect 406 4054 407 4058
rect 367 4004 407 4054
rect 367 4000 378 4004
rect 382 4000 390 4004
rect 394 4000 402 4004
rect 406 4000 407 4004
rect 367 3998 407 4000
rect 367 3994 378 3998
rect 382 3994 390 3998
rect 394 3994 402 3998
rect 406 3994 407 3998
rect 367 3992 407 3994
rect 367 3988 378 3992
rect 382 3988 390 3992
rect 394 3988 402 3992
rect 406 3988 407 3992
rect 367 3986 407 3988
rect 367 3982 378 3986
rect 382 3982 390 3986
rect 394 3982 402 3986
rect 406 3982 407 3986
rect 367 3980 407 3982
rect 367 3976 378 3980
rect 382 3976 390 3980
rect 394 3976 402 3980
rect 406 3976 407 3980
rect 367 3974 407 3976
rect 367 3970 378 3974
rect 382 3970 390 3974
rect 394 3970 402 3974
rect 406 3970 407 3974
rect 367 3968 407 3970
rect 367 3964 390 3968
rect 394 3964 402 3968
rect 406 3964 407 3968
rect 367 3620 407 3964
rect 367 3616 390 3620
rect 394 3616 402 3620
rect 406 3616 407 3620
rect 367 3614 407 3616
rect 367 3610 378 3614
rect 382 3610 390 3614
rect 394 3610 402 3614
rect 406 3610 407 3614
rect 367 3608 407 3610
rect 367 3604 378 3608
rect 382 3604 390 3608
rect 394 3604 402 3608
rect 406 3604 407 3608
rect 367 3602 407 3604
rect 367 3598 378 3602
rect 382 3598 390 3602
rect 394 3598 402 3602
rect 406 3598 407 3602
rect 367 3596 407 3598
rect 367 3592 378 3596
rect 382 3592 390 3596
rect 394 3592 402 3596
rect 406 3592 407 3596
rect 367 3590 407 3592
rect 367 3586 378 3590
rect 382 3586 390 3590
rect 394 3586 402 3590
rect 406 3586 407 3590
rect 367 3584 407 3586
rect 367 3580 378 3584
rect 382 3580 390 3584
rect 394 3580 402 3584
rect 406 3580 407 3584
rect 367 3530 407 3580
rect 367 3526 378 3530
rect 382 3526 390 3530
rect 394 3526 402 3530
rect 406 3526 407 3530
rect 367 3524 407 3526
rect 367 3520 378 3524
rect 382 3520 390 3524
rect 394 3520 402 3524
rect 406 3520 407 3524
rect 367 3518 407 3520
rect 367 3514 378 3518
rect 382 3514 390 3518
rect 394 3514 402 3518
rect 406 3514 407 3518
rect 367 3512 407 3514
rect 367 3508 378 3512
rect 382 3508 390 3512
rect 394 3508 402 3512
rect 406 3508 407 3512
rect 367 3506 407 3508
rect 367 3502 378 3506
rect 382 3502 390 3506
rect 394 3502 402 3506
rect 406 3502 407 3506
rect 367 3500 407 3502
rect 367 3496 378 3500
rect 382 3496 390 3500
rect 394 3496 402 3500
rect 406 3496 407 3500
rect 367 3494 407 3496
rect 367 3490 390 3494
rect 394 3490 402 3494
rect 406 3490 407 3494
rect 367 3146 407 3490
rect 367 3142 390 3146
rect 394 3142 402 3146
rect 406 3142 407 3146
rect 367 3140 407 3142
rect 367 3136 378 3140
rect 382 3136 390 3140
rect 394 3136 402 3140
rect 406 3136 407 3140
rect 367 3134 407 3136
rect 367 3130 378 3134
rect 382 3130 390 3134
rect 394 3130 402 3134
rect 406 3130 407 3134
rect 367 3128 407 3130
rect 367 3124 378 3128
rect 382 3124 390 3128
rect 394 3124 402 3128
rect 406 3124 407 3128
rect 367 3122 407 3124
rect 367 3118 378 3122
rect 382 3118 390 3122
rect 394 3118 402 3122
rect 406 3118 407 3122
rect 367 3116 407 3118
rect 367 3112 378 3116
rect 382 3112 390 3116
rect 394 3112 402 3116
rect 406 3112 407 3116
rect 367 3110 407 3112
rect 367 3106 378 3110
rect 382 3106 390 3110
rect 394 3106 402 3110
rect 406 3106 407 3110
rect 367 3056 407 3106
rect 367 3052 378 3056
rect 382 3052 390 3056
rect 394 3052 402 3056
rect 406 3052 407 3056
rect 367 3050 407 3052
rect 367 3046 378 3050
rect 382 3046 390 3050
rect 394 3046 402 3050
rect 406 3046 407 3050
rect 367 3044 407 3046
rect 367 3040 378 3044
rect 382 3040 390 3044
rect 394 3040 402 3044
rect 406 3040 407 3044
rect 367 3038 407 3040
rect 367 3034 378 3038
rect 382 3034 390 3038
rect 394 3034 402 3038
rect 406 3034 407 3038
rect 367 3032 407 3034
rect 367 3028 378 3032
rect 382 3028 390 3032
rect 394 3028 402 3032
rect 406 3028 407 3032
rect 367 3026 407 3028
rect 367 3022 378 3026
rect 382 3022 390 3026
rect 394 3022 402 3026
rect 406 3022 407 3026
rect 367 3020 407 3022
rect 367 3016 390 3020
rect 394 3016 402 3020
rect 406 3016 407 3020
rect 367 2672 407 3016
rect 367 2668 390 2672
rect 394 2668 402 2672
rect 406 2668 407 2672
rect 367 2666 407 2668
rect 367 2662 378 2666
rect 382 2662 390 2666
rect 394 2662 402 2666
rect 406 2662 407 2666
rect 367 2660 407 2662
rect 367 2656 378 2660
rect 382 2656 390 2660
rect 394 2656 402 2660
rect 406 2656 407 2660
rect 367 2654 407 2656
rect 367 2650 378 2654
rect 382 2650 390 2654
rect 394 2650 402 2654
rect 406 2650 407 2654
rect 367 2648 407 2650
rect 367 2644 378 2648
rect 382 2644 390 2648
rect 394 2644 402 2648
rect 406 2644 407 2648
rect 367 2642 407 2644
rect 367 2638 378 2642
rect 382 2638 390 2642
rect 394 2638 402 2642
rect 406 2638 407 2642
rect 367 2636 407 2638
rect 367 2632 378 2636
rect 382 2632 390 2636
rect 394 2632 402 2636
rect 406 2632 407 2636
rect 367 2582 407 2632
rect 367 2578 378 2582
rect 382 2578 390 2582
rect 394 2578 402 2582
rect 406 2578 407 2582
rect 367 2576 407 2578
rect 367 2572 378 2576
rect 382 2572 390 2576
rect 394 2572 402 2576
rect 406 2572 407 2576
rect 367 2570 407 2572
rect 367 2566 378 2570
rect 382 2566 390 2570
rect 394 2566 402 2570
rect 406 2566 407 2570
rect 367 2564 407 2566
rect 367 2560 378 2564
rect 382 2560 390 2564
rect 394 2560 402 2564
rect 406 2560 407 2564
rect 367 2558 407 2560
rect 367 2554 378 2558
rect 382 2554 390 2558
rect 394 2554 402 2558
rect 406 2554 407 2558
rect 367 2552 407 2554
rect 367 2548 378 2552
rect 382 2548 390 2552
rect 394 2548 402 2552
rect 406 2548 407 2552
rect 367 2546 407 2548
rect 367 2542 390 2546
rect 394 2542 402 2546
rect 406 2542 407 2546
rect 367 2198 407 2542
rect 367 2194 390 2198
rect 394 2194 402 2198
rect 406 2194 407 2198
rect 367 2192 407 2194
rect 367 2188 378 2192
rect 382 2188 390 2192
rect 394 2188 402 2192
rect 406 2188 407 2192
rect 367 2186 407 2188
rect 367 2182 378 2186
rect 382 2182 390 2186
rect 394 2182 402 2186
rect 406 2182 407 2186
rect 367 2180 407 2182
rect 367 2176 378 2180
rect 382 2176 390 2180
rect 394 2176 402 2180
rect 406 2176 407 2180
rect 367 2174 407 2176
rect 367 2170 378 2174
rect 382 2170 390 2174
rect 394 2170 402 2174
rect 406 2170 407 2174
rect 367 2168 407 2170
rect 367 2164 378 2168
rect 382 2164 390 2168
rect 394 2164 402 2168
rect 406 2164 407 2168
rect 367 2162 407 2164
rect 367 2158 378 2162
rect 382 2158 390 2162
rect 394 2158 402 2162
rect 406 2158 407 2162
rect 367 2108 407 2158
rect 367 2104 378 2108
rect 382 2104 390 2108
rect 394 2104 402 2108
rect 406 2104 407 2108
rect 367 2102 407 2104
rect 367 2098 378 2102
rect 382 2098 390 2102
rect 394 2098 402 2102
rect 406 2098 407 2102
rect 367 2096 407 2098
rect 367 2092 378 2096
rect 382 2092 390 2096
rect 394 2092 402 2096
rect 406 2092 407 2096
rect 367 2090 407 2092
rect 367 2086 378 2090
rect 382 2086 390 2090
rect 394 2086 402 2090
rect 406 2086 407 2090
rect 367 2084 407 2086
rect 367 2080 378 2084
rect 382 2080 390 2084
rect 394 2080 402 2084
rect 406 2080 407 2084
rect 367 2078 407 2080
rect 367 2074 378 2078
rect 382 2074 390 2078
rect 394 2074 402 2078
rect 406 2074 407 2078
rect 367 2072 407 2074
rect 367 2068 390 2072
rect 394 2068 402 2072
rect 406 2068 407 2072
rect 367 1724 407 2068
rect 367 1720 390 1724
rect 394 1720 402 1724
rect 406 1720 407 1724
rect 367 1718 407 1720
rect 367 1714 378 1718
rect 382 1714 390 1718
rect 394 1714 402 1718
rect 406 1714 407 1718
rect 367 1712 407 1714
rect 367 1708 378 1712
rect 382 1708 390 1712
rect 394 1708 402 1712
rect 406 1708 407 1712
rect 367 1706 407 1708
rect 367 1702 378 1706
rect 382 1702 390 1706
rect 394 1702 402 1706
rect 406 1702 407 1706
rect 367 1700 407 1702
rect 367 1696 378 1700
rect 382 1696 390 1700
rect 394 1696 402 1700
rect 406 1696 407 1700
rect 367 1694 407 1696
rect 367 1690 378 1694
rect 382 1690 390 1694
rect 394 1690 402 1694
rect 406 1690 407 1694
rect 367 1688 407 1690
rect 367 1684 378 1688
rect 382 1684 390 1688
rect 394 1684 402 1688
rect 406 1684 407 1688
rect 367 1634 407 1684
rect 367 1630 378 1634
rect 382 1630 390 1634
rect 394 1630 402 1634
rect 406 1630 407 1634
rect 367 1628 407 1630
rect 367 1624 378 1628
rect 382 1624 390 1628
rect 394 1624 402 1628
rect 406 1624 407 1628
rect 367 1622 407 1624
rect 367 1618 378 1622
rect 382 1618 390 1622
rect 394 1618 402 1622
rect 406 1618 407 1622
rect 367 1616 407 1618
rect 367 1612 378 1616
rect 382 1612 390 1616
rect 394 1612 402 1616
rect 406 1612 407 1616
rect 367 1610 407 1612
rect 367 1606 378 1610
rect 382 1606 390 1610
rect 394 1606 402 1610
rect 406 1606 407 1610
rect 367 1604 407 1606
rect 367 1600 378 1604
rect 382 1600 390 1604
rect 394 1600 402 1604
rect 406 1600 407 1604
rect 367 1598 407 1600
rect 367 1594 390 1598
rect 394 1594 402 1598
rect 406 1594 407 1598
rect 367 1250 407 1594
rect 367 1246 390 1250
rect 394 1246 402 1250
rect 406 1246 407 1250
rect 367 1244 407 1246
rect 367 1240 378 1244
rect 382 1240 390 1244
rect 394 1240 402 1244
rect 406 1240 407 1244
rect 367 1238 407 1240
rect 367 1234 378 1238
rect 382 1234 390 1238
rect 394 1234 402 1238
rect 406 1234 407 1238
rect 367 1232 407 1234
rect 367 1228 378 1232
rect 382 1228 390 1232
rect 394 1228 402 1232
rect 406 1228 407 1232
rect 367 1226 407 1228
rect 367 1222 378 1226
rect 382 1222 390 1226
rect 394 1222 402 1226
rect 406 1222 407 1226
rect 367 1220 407 1222
rect 367 1216 378 1220
rect 382 1216 390 1220
rect 394 1216 402 1220
rect 406 1216 407 1220
rect 367 1214 407 1216
rect 367 1210 378 1214
rect 382 1210 390 1214
rect 394 1210 402 1214
rect 406 1210 407 1214
rect 367 1160 407 1210
rect 367 1156 378 1160
rect 382 1156 390 1160
rect 394 1156 402 1160
rect 406 1156 407 1160
rect 367 1154 407 1156
rect 367 1150 378 1154
rect 382 1150 390 1154
rect 394 1150 402 1154
rect 406 1150 407 1154
rect 367 1148 407 1150
rect 367 1144 378 1148
rect 382 1144 390 1148
rect 394 1144 402 1148
rect 406 1144 407 1148
rect 367 1142 407 1144
rect 367 1138 378 1142
rect 382 1138 390 1142
rect 394 1138 402 1142
rect 406 1138 407 1142
rect 367 1136 407 1138
rect 367 1132 378 1136
rect 382 1132 390 1136
rect 394 1132 402 1136
rect 406 1132 407 1136
rect 367 1130 407 1132
rect 367 1126 378 1130
rect 382 1126 390 1130
rect 394 1126 402 1130
rect 406 1126 407 1130
rect 367 1124 407 1126
rect 367 1120 390 1124
rect 394 1120 402 1124
rect 406 1120 407 1124
rect 367 776 407 1120
rect 367 772 390 776
rect 394 772 402 776
rect 406 772 407 776
rect 367 770 407 772
rect 367 766 378 770
rect 382 766 390 770
rect 394 766 402 770
rect 406 766 407 770
rect 367 764 407 766
rect 367 760 378 764
rect 382 760 390 764
rect 394 760 402 764
rect 406 760 407 764
rect 367 758 407 760
rect 367 754 378 758
rect 382 754 390 758
rect 394 754 402 758
rect 406 754 407 758
rect 367 752 407 754
rect 367 748 378 752
rect 382 748 390 752
rect 394 748 402 752
rect 406 748 407 752
rect 367 746 407 748
rect 367 742 378 746
rect 382 742 390 746
rect 394 742 402 746
rect 406 742 407 746
rect 367 740 407 742
rect 367 736 378 740
rect 382 736 390 740
rect 394 736 402 740
rect 406 736 407 740
rect 367 686 407 736
rect 367 682 378 686
rect 382 682 390 686
rect 394 682 402 686
rect 406 682 407 686
rect 367 680 407 682
rect 367 676 378 680
rect 382 676 390 680
rect 394 676 402 680
rect 406 676 407 680
rect 367 674 407 676
rect 367 670 378 674
rect 382 670 390 674
rect 394 670 402 674
rect 406 670 407 674
rect 367 668 407 670
rect 367 664 378 668
rect 382 664 390 668
rect 394 664 402 668
rect 406 664 407 668
rect 367 662 407 664
rect 367 658 378 662
rect 382 658 390 662
rect 394 658 402 662
rect 406 658 407 662
rect 367 656 407 658
rect 367 652 378 656
rect 382 652 390 656
rect 394 652 402 656
rect 406 652 407 656
rect 367 650 407 652
rect 367 646 390 650
rect 394 646 402 650
rect 406 646 407 650
rect 367 302 407 646
rect 367 298 390 302
rect 394 298 402 302
rect 406 298 407 302
rect 367 296 407 298
rect 367 292 378 296
rect 382 292 390 296
rect 394 292 402 296
rect 406 292 407 296
rect 367 290 407 292
rect 367 286 378 290
rect 382 286 390 290
rect 394 286 402 290
rect 406 286 407 290
rect 367 284 407 286
rect 367 280 378 284
rect 382 280 390 284
rect 394 280 402 284
rect 406 280 407 284
rect 367 278 407 280
rect 367 274 378 278
rect 382 274 390 278
rect 394 274 402 278
rect 406 274 407 278
rect 367 272 407 274
rect 367 268 378 272
rect 382 268 390 272
rect 394 268 402 272
rect 406 268 407 272
rect 367 266 407 268
rect 367 262 378 266
rect 382 262 390 266
rect 394 262 402 266
rect 406 262 407 266
rect 367 212 407 262
rect 367 208 378 212
rect 382 208 390 212
rect 394 208 402 212
rect 406 208 407 212
rect 367 206 407 208
rect 367 202 378 206
rect 382 202 390 206
rect 394 202 402 206
rect 406 202 407 206
rect 367 200 407 202
rect 367 196 378 200
rect 382 196 390 200
rect 394 196 402 200
rect 406 196 407 200
rect 367 194 407 196
rect 367 190 378 194
rect 382 190 390 194
rect 394 190 402 194
rect 406 190 407 194
rect 367 188 407 190
rect 367 184 378 188
rect 382 184 390 188
rect 394 184 402 188
rect 406 184 407 188
rect 367 182 407 184
rect 367 178 378 182
rect 382 178 390 182
rect 394 178 402 182
rect 406 178 407 182
rect 367 176 407 178
rect 367 172 390 176
rect 394 172 402 176
rect 406 172 407 176
rect 367 40 407 172
rect 411 4180 451 4182
rect 411 4146 413 4180
rect 447 4146 451 4180
rect 411 4138 451 4146
rect 411 4134 412 4138
rect 421 4134 423 4138
rect 427 4134 429 4138
rect 433 4134 435 4138
rect 439 4134 441 4138
rect 450 4134 451 4138
rect 411 4132 451 4134
rect 411 4128 412 4132
rect 421 4128 423 4132
rect 427 4128 429 4132
rect 433 4128 435 4132
rect 439 4128 441 4132
rect 450 4128 451 4132
rect 411 4126 451 4128
rect 411 4122 412 4126
rect 421 4122 423 4126
rect 427 4122 429 4126
rect 433 4122 435 4126
rect 439 4122 441 4126
rect 450 4122 451 4126
rect 411 4120 451 4122
rect 411 4116 412 4120
rect 421 4116 423 4120
rect 427 4116 429 4120
rect 433 4116 435 4120
rect 439 4116 441 4120
rect 450 4116 451 4120
rect 411 4114 451 4116
rect 411 4110 412 4114
rect 421 4110 423 4114
rect 427 4110 429 4114
rect 433 4110 435 4114
rect 439 4110 441 4114
rect 450 4110 451 4114
rect 411 4108 451 4110
rect 411 4104 412 4108
rect 421 4104 423 4108
rect 427 4104 429 4108
rect 433 4104 435 4108
rect 439 4104 441 4108
rect 450 4104 451 4108
rect 411 4102 451 4104
rect 411 4098 412 4102
rect 421 4098 423 4102
rect 427 4098 429 4102
rect 433 4098 435 4102
rect 439 4098 441 4102
rect 450 4098 451 4102
rect 411 3960 451 4098
rect 411 3956 412 3960
rect 421 3956 423 3960
rect 427 3956 429 3960
rect 433 3956 435 3960
rect 439 3956 441 3960
rect 450 3956 451 3960
rect 411 3954 451 3956
rect 411 3950 412 3954
rect 421 3950 423 3954
rect 427 3950 429 3954
rect 433 3950 435 3954
rect 439 3950 441 3954
rect 450 3950 451 3954
rect 411 3948 451 3950
rect 411 3944 412 3948
rect 421 3944 423 3948
rect 427 3944 429 3948
rect 433 3944 435 3948
rect 439 3944 441 3948
rect 450 3944 451 3948
rect 411 3942 451 3944
rect 411 3938 412 3942
rect 421 3938 423 3942
rect 427 3938 429 3942
rect 433 3938 435 3942
rect 439 3938 441 3942
rect 450 3938 451 3942
rect 411 3936 451 3938
rect 411 3932 412 3936
rect 421 3932 423 3936
rect 427 3932 429 3936
rect 433 3932 435 3936
rect 439 3932 441 3936
rect 450 3932 451 3936
rect 411 3930 451 3932
rect 411 3926 412 3930
rect 421 3926 423 3930
rect 427 3926 429 3930
rect 433 3926 435 3930
rect 439 3926 441 3930
rect 450 3926 451 3930
rect 411 3924 451 3926
rect 411 3920 412 3924
rect 421 3920 423 3924
rect 427 3920 429 3924
rect 433 3920 435 3924
rect 439 3920 441 3924
rect 450 3920 451 3924
rect 411 3664 451 3920
rect 411 3660 412 3664
rect 421 3660 423 3664
rect 427 3660 429 3664
rect 433 3660 435 3664
rect 439 3660 441 3664
rect 450 3660 451 3664
rect 411 3658 451 3660
rect 411 3654 412 3658
rect 421 3654 423 3658
rect 427 3654 429 3658
rect 433 3654 435 3658
rect 439 3654 441 3658
rect 450 3654 451 3658
rect 411 3652 451 3654
rect 411 3648 412 3652
rect 421 3648 423 3652
rect 427 3648 429 3652
rect 433 3648 435 3652
rect 439 3648 441 3652
rect 450 3648 451 3652
rect 411 3646 451 3648
rect 411 3642 412 3646
rect 421 3642 423 3646
rect 427 3642 429 3646
rect 433 3642 435 3646
rect 439 3642 441 3646
rect 450 3642 451 3646
rect 411 3640 451 3642
rect 411 3636 412 3640
rect 421 3636 423 3640
rect 427 3636 429 3640
rect 433 3636 435 3640
rect 439 3636 441 3640
rect 450 3636 451 3640
rect 411 3634 451 3636
rect 411 3630 412 3634
rect 421 3630 423 3634
rect 427 3630 429 3634
rect 433 3630 435 3634
rect 439 3630 441 3634
rect 450 3630 451 3634
rect 411 3628 451 3630
rect 411 3624 412 3628
rect 421 3624 423 3628
rect 427 3624 429 3628
rect 433 3624 435 3628
rect 439 3624 441 3628
rect 450 3624 451 3628
rect 411 3486 451 3624
rect 411 3482 412 3486
rect 421 3482 423 3486
rect 427 3482 429 3486
rect 433 3482 435 3486
rect 439 3482 441 3486
rect 450 3482 451 3486
rect 411 3480 451 3482
rect 411 3476 412 3480
rect 421 3476 423 3480
rect 427 3476 429 3480
rect 433 3476 435 3480
rect 439 3476 441 3480
rect 450 3476 451 3480
rect 411 3474 451 3476
rect 411 3470 412 3474
rect 421 3470 423 3474
rect 427 3470 429 3474
rect 433 3470 435 3474
rect 439 3470 441 3474
rect 450 3470 451 3474
rect 411 3468 451 3470
rect 411 3464 412 3468
rect 421 3464 423 3468
rect 427 3464 429 3468
rect 433 3464 435 3468
rect 439 3464 441 3468
rect 450 3464 451 3468
rect 411 3462 451 3464
rect 411 3458 412 3462
rect 421 3458 423 3462
rect 427 3458 429 3462
rect 433 3458 435 3462
rect 439 3458 441 3462
rect 450 3458 451 3462
rect 411 3456 451 3458
rect 411 3452 412 3456
rect 421 3452 423 3456
rect 427 3452 429 3456
rect 433 3452 435 3456
rect 439 3452 441 3456
rect 450 3452 451 3456
rect 411 3450 451 3452
rect 411 3446 412 3450
rect 421 3446 423 3450
rect 427 3446 429 3450
rect 433 3446 435 3450
rect 439 3446 441 3450
rect 450 3446 451 3450
rect 411 3190 451 3446
rect 411 3186 412 3190
rect 421 3186 423 3190
rect 427 3186 429 3190
rect 433 3186 435 3190
rect 439 3186 441 3190
rect 450 3186 451 3190
rect 411 3184 451 3186
rect 411 3180 412 3184
rect 421 3180 423 3184
rect 427 3180 429 3184
rect 433 3180 435 3184
rect 439 3180 441 3184
rect 450 3180 451 3184
rect 411 3178 451 3180
rect 411 3174 412 3178
rect 421 3174 423 3178
rect 427 3174 429 3178
rect 433 3174 435 3178
rect 439 3174 441 3178
rect 450 3174 451 3178
rect 411 3172 451 3174
rect 411 3168 412 3172
rect 421 3168 423 3172
rect 427 3168 429 3172
rect 433 3168 435 3172
rect 439 3168 441 3172
rect 450 3168 451 3172
rect 411 3166 451 3168
rect 411 3162 412 3166
rect 421 3162 423 3166
rect 427 3162 429 3166
rect 433 3162 435 3166
rect 439 3162 441 3166
rect 450 3162 451 3166
rect 411 3160 451 3162
rect 411 3156 412 3160
rect 421 3156 423 3160
rect 427 3156 429 3160
rect 433 3156 435 3160
rect 439 3156 441 3160
rect 450 3156 451 3160
rect 411 3154 451 3156
rect 411 3150 412 3154
rect 421 3150 423 3154
rect 427 3150 429 3154
rect 433 3150 435 3154
rect 439 3150 441 3154
rect 450 3150 451 3154
rect 411 3012 451 3150
rect 411 3008 412 3012
rect 421 3008 423 3012
rect 427 3008 429 3012
rect 433 3008 435 3012
rect 439 3008 441 3012
rect 450 3008 451 3012
rect 411 3006 451 3008
rect 411 3002 412 3006
rect 421 3002 423 3006
rect 427 3002 429 3006
rect 433 3002 435 3006
rect 439 3002 441 3006
rect 450 3002 451 3006
rect 411 3000 451 3002
rect 411 2996 412 3000
rect 421 2996 423 3000
rect 427 2996 429 3000
rect 433 2996 435 3000
rect 439 2996 441 3000
rect 450 2996 451 3000
rect 411 2994 451 2996
rect 411 2990 412 2994
rect 421 2990 423 2994
rect 427 2990 429 2994
rect 433 2990 435 2994
rect 439 2990 441 2994
rect 450 2990 451 2994
rect 411 2988 451 2990
rect 411 2984 412 2988
rect 421 2984 423 2988
rect 427 2984 429 2988
rect 433 2984 435 2988
rect 439 2984 441 2988
rect 450 2984 451 2988
rect 411 2982 451 2984
rect 411 2978 412 2982
rect 421 2978 423 2982
rect 427 2978 429 2982
rect 433 2978 435 2982
rect 439 2978 441 2982
rect 450 2978 451 2982
rect 411 2976 451 2978
rect 411 2972 412 2976
rect 421 2972 423 2976
rect 427 2972 429 2976
rect 433 2972 435 2976
rect 439 2972 441 2976
rect 450 2972 451 2976
rect 411 2716 451 2972
rect 411 2712 412 2716
rect 421 2712 423 2716
rect 427 2712 429 2716
rect 433 2712 435 2716
rect 439 2712 441 2716
rect 450 2712 451 2716
rect 411 2710 451 2712
rect 411 2706 412 2710
rect 421 2706 423 2710
rect 427 2706 429 2710
rect 433 2706 435 2710
rect 439 2706 441 2710
rect 450 2706 451 2710
rect 411 2704 451 2706
rect 411 2700 412 2704
rect 421 2700 423 2704
rect 427 2700 429 2704
rect 433 2700 435 2704
rect 439 2700 441 2704
rect 450 2700 451 2704
rect 411 2698 451 2700
rect 411 2694 412 2698
rect 421 2694 423 2698
rect 427 2694 429 2698
rect 433 2694 435 2698
rect 439 2694 441 2698
rect 450 2694 451 2698
rect 411 2692 451 2694
rect 411 2688 412 2692
rect 421 2688 423 2692
rect 427 2688 429 2692
rect 433 2688 435 2692
rect 439 2688 441 2692
rect 450 2688 451 2692
rect 411 2686 451 2688
rect 411 2682 412 2686
rect 421 2682 423 2686
rect 427 2682 429 2686
rect 433 2682 435 2686
rect 439 2682 441 2686
rect 450 2682 451 2686
rect 411 2680 451 2682
rect 411 2676 412 2680
rect 421 2676 423 2680
rect 427 2676 429 2680
rect 433 2676 435 2680
rect 439 2676 441 2680
rect 450 2676 451 2680
rect 411 2538 451 2676
rect 411 2534 412 2538
rect 421 2534 423 2538
rect 427 2534 429 2538
rect 433 2534 435 2538
rect 439 2534 441 2538
rect 450 2534 451 2538
rect 411 2532 451 2534
rect 411 2528 412 2532
rect 421 2528 423 2532
rect 427 2528 429 2532
rect 433 2528 435 2532
rect 439 2528 441 2532
rect 450 2528 451 2532
rect 411 2526 451 2528
rect 411 2522 412 2526
rect 421 2522 423 2526
rect 427 2522 429 2526
rect 433 2522 435 2526
rect 439 2522 441 2526
rect 450 2522 451 2526
rect 411 2520 451 2522
rect 411 2516 412 2520
rect 421 2516 423 2520
rect 427 2516 429 2520
rect 433 2516 435 2520
rect 439 2516 441 2520
rect 450 2516 451 2520
rect 411 2514 451 2516
rect 411 2510 412 2514
rect 421 2510 423 2514
rect 427 2510 429 2514
rect 433 2510 435 2514
rect 439 2510 441 2514
rect 450 2510 451 2514
rect 411 2508 451 2510
rect 411 2504 412 2508
rect 421 2504 423 2508
rect 427 2504 429 2508
rect 433 2504 435 2508
rect 439 2504 441 2508
rect 450 2504 451 2508
rect 411 2502 451 2504
rect 411 2498 412 2502
rect 421 2498 423 2502
rect 427 2498 429 2502
rect 433 2498 435 2502
rect 439 2498 441 2502
rect 450 2498 451 2502
rect 411 2242 451 2498
rect 411 2238 412 2242
rect 421 2238 423 2242
rect 427 2238 429 2242
rect 433 2238 435 2242
rect 439 2238 441 2242
rect 450 2238 451 2242
rect 411 2236 451 2238
rect 411 2232 412 2236
rect 421 2232 423 2236
rect 427 2232 429 2236
rect 433 2232 435 2236
rect 439 2232 441 2236
rect 450 2232 451 2236
rect 411 2230 451 2232
rect 411 2226 412 2230
rect 421 2226 423 2230
rect 427 2226 429 2230
rect 433 2226 435 2230
rect 439 2226 441 2230
rect 450 2226 451 2230
rect 411 2224 451 2226
rect 411 2220 412 2224
rect 421 2220 423 2224
rect 427 2220 429 2224
rect 433 2220 435 2224
rect 439 2220 441 2224
rect 450 2220 451 2224
rect 411 2218 451 2220
rect 411 2214 412 2218
rect 421 2214 423 2218
rect 427 2214 429 2218
rect 433 2214 435 2218
rect 439 2214 441 2218
rect 450 2214 451 2218
rect 411 2212 451 2214
rect 411 2208 412 2212
rect 421 2208 423 2212
rect 427 2208 429 2212
rect 433 2208 435 2212
rect 439 2208 441 2212
rect 450 2208 451 2212
rect 411 2206 451 2208
rect 411 2202 412 2206
rect 421 2202 423 2206
rect 427 2202 429 2206
rect 433 2202 435 2206
rect 439 2202 441 2206
rect 450 2202 451 2206
rect 411 2064 451 2202
rect 411 2060 412 2064
rect 421 2060 423 2064
rect 427 2060 429 2064
rect 433 2060 435 2064
rect 439 2060 441 2064
rect 450 2060 451 2064
rect 411 2058 451 2060
rect 411 2054 412 2058
rect 421 2054 423 2058
rect 427 2054 429 2058
rect 433 2054 435 2058
rect 439 2054 441 2058
rect 450 2054 451 2058
rect 411 2052 451 2054
rect 411 2048 412 2052
rect 421 2048 423 2052
rect 427 2048 429 2052
rect 433 2048 435 2052
rect 439 2048 441 2052
rect 450 2048 451 2052
rect 411 2046 451 2048
rect 411 2042 412 2046
rect 421 2042 423 2046
rect 427 2042 429 2046
rect 433 2042 435 2046
rect 439 2042 441 2046
rect 450 2042 451 2046
rect 411 2040 451 2042
rect 411 2036 412 2040
rect 421 2036 423 2040
rect 427 2036 429 2040
rect 433 2036 435 2040
rect 439 2036 441 2040
rect 450 2036 451 2040
rect 411 2034 451 2036
rect 411 2030 412 2034
rect 421 2030 423 2034
rect 427 2030 429 2034
rect 433 2030 435 2034
rect 439 2030 441 2034
rect 450 2030 451 2034
rect 411 2028 451 2030
rect 411 2024 412 2028
rect 421 2024 423 2028
rect 427 2024 429 2028
rect 433 2024 435 2028
rect 439 2024 441 2028
rect 450 2024 451 2028
rect 411 1768 451 2024
rect 411 1764 412 1768
rect 421 1764 423 1768
rect 427 1764 429 1768
rect 433 1764 435 1768
rect 439 1764 441 1768
rect 450 1764 451 1768
rect 411 1762 451 1764
rect 411 1758 412 1762
rect 421 1758 423 1762
rect 427 1758 429 1762
rect 433 1758 435 1762
rect 439 1758 441 1762
rect 450 1758 451 1762
rect 411 1756 451 1758
rect 411 1752 412 1756
rect 421 1752 423 1756
rect 427 1752 429 1756
rect 433 1752 435 1756
rect 439 1752 441 1756
rect 450 1752 451 1756
rect 411 1750 451 1752
rect 411 1746 412 1750
rect 421 1746 423 1750
rect 427 1746 429 1750
rect 433 1746 435 1750
rect 439 1746 441 1750
rect 450 1746 451 1750
rect 411 1744 451 1746
rect 411 1740 412 1744
rect 421 1740 423 1744
rect 427 1740 429 1744
rect 433 1740 435 1744
rect 439 1740 441 1744
rect 450 1740 451 1744
rect 411 1738 451 1740
rect 411 1734 412 1738
rect 421 1734 423 1738
rect 427 1734 429 1738
rect 433 1734 435 1738
rect 439 1734 441 1738
rect 450 1734 451 1738
rect 411 1732 451 1734
rect 411 1728 412 1732
rect 421 1728 423 1732
rect 427 1728 429 1732
rect 433 1728 435 1732
rect 439 1728 441 1732
rect 450 1728 451 1732
rect 411 1590 451 1728
rect 411 1586 412 1590
rect 421 1586 423 1590
rect 427 1586 429 1590
rect 433 1586 435 1590
rect 439 1586 441 1590
rect 450 1586 451 1590
rect 411 1584 451 1586
rect 411 1580 412 1584
rect 421 1580 423 1584
rect 427 1580 429 1584
rect 433 1580 435 1584
rect 439 1580 441 1584
rect 450 1580 451 1584
rect 411 1578 451 1580
rect 411 1574 412 1578
rect 421 1574 423 1578
rect 427 1574 429 1578
rect 433 1574 435 1578
rect 439 1574 441 1578
rect 450 1574 451 1578
rect 411 1572 451 1574
rect 411 1568 412 1572
rect 421 1568 423 1572
rect 427 1568 429 1572
rect 433 1568 435 1572
rect 439 1568 441 1572
rect 450 1568 451 1572
rect 411 1566 451 1568
rect 411 1562 412 1566
rect 421 1562 423 1566
rect 427 1562 429 1566
rect 433 1562 435 1566
rect 439 1562 441 1566
rect 450 1562 451 1566
rect 411 1560 451 1562
rect 411 1556 412 1560
rect 421 1556 423 1560
rect 427 1556 429 1560
rect 433 1556 435 1560
rect 439 1556 441 1560
rect 450 1556 451 1560
rect 411 1554 451 1556
rect 411 1550 412 1554
rect 421 1550 423 1554
rect 427 1550 429 1554
rect 433 1550 435 1554
rect 439 1550 441 1554
rect 450 1550 451 1554
rect 411 1294 451 1550
rect 411 1290 412 1294
rect 421 1290 423 1294
rect 427 1290 429 1294
rect 433 1290 435 1294
rect 439 1290 441 1294
rect 450 1290 451 1294
rect 411 1288 451 1290
rect 411 1284 412 1288
rect 421 1284 423 1288
rect 427 1284 429 1288
rect 433 1284 435 1288
rect 439 1284 441 1288
rect 450 1284 451 1288
rect 411 1282 451 1284
rect 411 1278 412 1282
rect 421 1278 423 1282
rect 427 1278 429 1282
rect 433 1278 435 1282
rect 439 1278 441 1282
rect 450 1278 451 1282
rect 411 1276 451 1278
rect 411 1272 412 1276
rect 421 1272 423 1276
rect 427 1272 429 1276
rect 433 1272 435 1276
rect 439 1272 441 1276
rect 450 1272 451 1276
rect 411 1270 451 1272
rect 411 1266 412 1270
rect 421 1266 423 1270
rect 427 1266 429 1270
rect 433 1266 435 1270
rect 439 1266 441 1270
rect 450 1266 451 1270
rect 411 1264 451 1266
rect 411 1260 412 1264
rect 421 1260 423 1264
rect 427 1260 429 1264
rect 433 1260 435 1264
rect 439 1260 441 1264
rect 450 1260 451 1264
rect 411 1258 451 1260
rect 411 1254 412 1258
rect 421 1254 423 1258
rect 427 1254 429 1258
rect 433 1254 435 1258
rect 439 1254 441 1258
rect 450 1254 451 1258
rect 411 1116 451 1254
rect 411 1112 412 1116
rect 421 1112 423 1116
rect 427 1112 429 1116
rect 433 1112 435 1116
rect 439 1112 441 1116
rect 450 1112 451 1116
rect 411 1110 451 1112
rect 411 1106 412 1110
rect 421 1106 423 1110
rect 427 1106 429 1110
rect 433 1106 435 1110
rect 439 1106 441 1110
rect 450 1106 451 1110
rect 411 1104 451 1106
rect 411 1100 412 1104
rect 421 1100 423 1104
rect 427 1100 429 1104
rect 433 1100 435 1104
rect 439 1100 441 1104
rect 450 1100 451 1104
rect 411 1098 451 1100
rect 411 1094 412 1098
rect 421 1094 423 1098
rect 427 1094 429 1098
rect 433 1094 435 1098
rect 439 1094 441 1098
rect 450 1094 451 1098
rect 411 1092 451 1094
rect 411 1088 412 1092
rect 421 1088 423 1092
rect 427 1088 429 1092
rect 433 1088 435 1092
rect 439 1088 441 1092
rect 450 1088 451 1092
rect 411 1086 451 1088
rect 411 1082 412 1086
rect 421 1082 423 1086
rect 427 1082 429 1086
rect 433 1082 435 1086
rect 439 1082 441 1086
rect 450 1082 451 1086
rect 411 1080 451 1082
rect 411 1076 412 1080
rect 421 1076 423 1080
rect 427 1076 429 1080
rect 433 1076 435 1080
rect 439 1076 441 1080
rect 450 1076 451 1080
rect 411 820 451 1076
rect 411 816 412 820
rect 421 816 423 820
rect 427 816 429 820
rect 433 816 435 820
rect 439 816 441 820
rect 450 816 451 820
rect 411 814 451 816
rect 411 810 412 814
rect 421 810 423 814
rect 427 810 429 814
rect 433 810 435 814
rect 439 810 441 814
rect 450 810 451 814
rect 411 808 451 810
rect 411 804 412 808
rect 421 804 423 808
rect 427 804 429 808
rect 433 804 435 808
rect 439 804 441 808
rect 450 804 451 808
rect 411 802 451 804
rect 411 798 412 802
rect 421 798 423 802
rect 427 798 429 802
rect 433 798 435 802
rect 439 798 441 802
rect 450 798 451 802
rect 411 796 451 798
rect 411 792 412 796
rect 421 792 423 796
rect 427 792 429 796
rect 433 792 435 796
rect 439 792 441 796
rect 450 792 451 796
rect 411 790 451 792
rect 411 786 412 790
rect 421 786 423 790
rect 427 786 429 790
rect 433 786 435 790
rect 439 786 441 790
rect 450 786 451 790
rect 411 784 451 786
rect 411 780 412 784
rect 421 780 423 784
rect 427 780 429 784
rect 433 780 435 784
rect 439 780 441 784
rect 450 780 451 784
rect 411 642 451 780
rect 411 638 412 642
rect 421 638 423 642
rect 427 638 429 642
rect 433 638 435 642
rect 439 638 441 642
rect 450 638 451 642
rect 411 636 451 638
rect 411 632 412 636
rect 421 632 423 636
rect 427 632 429 636
rect 433 632 435 636
rect 439 632 441 636
rect 450 632 451 636
rect 411 630 451 632
rect 411 626 412 630
rect 421 626 423 630
rect 427 626 429 630
rect 433 626 435 630
rect 439 626 441 630
rect 450 626 451 630
rect 411 624 451 626
rect 411 620 412 624
rect 421 620 423 624
rect 427 620 429 624
rect 433 620 435 624
rect 439 620 441 624
rect 450 620 451 624
rect 411 618 451 620
rect 411 614 412 618
rect 421 614 423 618
rect 427 614 429 618
rect 433 614 435 618
rect 439 614 441 618
rect 450 614 451 618
rect 411 612 451 614
rect 411 608 412 612
rect 421 608 423 612
rect 427 608 429 612
rect 433 608 435 612
rect 439 608 441 612
rect 450 608 451 612
rect 411 606 451 608
rect 411 602 412 606
rect 421 602 423 606
rect 427 602 429 606
rect 433 602 435 606
rect 439 602 441 606
rect 450 602 451 606
rect 411 346 451 602
rect 411 342 412 346
rect 421 342 423 346
rect 427 342 429 346
rect 433 342 435 346
rect 439 342 441 346
rect 450 342 451 346
rect 411 340 451 342
rect 411 336 412 340
rect 421 336 423 340
rect 427 336 429 340
rect 433 336 435 340
rect 439 336 441 340
rect 450 336 451 340
rect 411 334 451 336
rect 411 330 412 334
rect 421 330 423 334
rect 427 330 429 334
rect 433 330 435 334
rect 439 330 441 334
rect 450 330 451 334
rect 411 328 451 330
rect 411 324 412 328
rect 421 324 423 328
rect 427 324 429 328
rect 433 324 435 328
rect 439 324 441 328
rect 450 324 451 328
rect 411 322 451 324
rect 411 318 412 322
rect 421 318 423 322
rect 427 318 429 322
rect 433 318 435 322
rect 439 318 441 322
rect 450 318 451 322
rect 411 316 451 318
rect 411 312 412 316
rect 421 312 423 316
rect 427 312 429 316
rect 433 312 435 316
rect 439 312 441 316
rect 450 312 451 316
rect 411 310 451 312
rect 411 306 412 310
rect 421 306 423 310
rect 427 306 429 310
rect 433 306 435 310
rect 439 306 441 310
rect 450 306 451 310
rect 411 168 451 306
rect 411 164 412 168
rect 421 164 423 168
rect 427 164 429 168
rect 433 164 435 168
rect 439 164 441 168
rect 450 164 451 168
rect 411 162 451 164
rect 411 158 412 162
rect 421 158 423 162
rect 427 158 429 162
rect 433 158 435 162
rect 439 158 441 162
rect 450 158 451 162
rect 411 156 451 158
rect 411 152 412 156
rect 421 152 423 156
rect 427 152 429 156
rect 433 152 435 156
rect 439 152 441 156
rect 450 152 451 156
rect 411 150 451 152
rect 411 146 412 150
rect 421 146 423 150
rect 427 146 429 150
rect 433 146 435 150
rect 439 146 441 150
rect 450 146 451 150
rect 411 144 451 146
rect 411 140 412 144
rect 421 140 423 144
rect 427 140 429 144
rect 433 140 435 144
rect 439 140 441 144
rect 450 140 451 144
rect 411 138 451 140
rect 411 134 412 138
rect 421 134 423 138
rect 427 134 429 138
rect 433 134 435 138
rect 439 134 441 138
rect 450 134 451 138
rect 411 132 451 134
rect 411 128 412 132
rect 421 128 423 132
rect 427 128 429 132
rect 433 128 435 132
rect 439 128 441 132
rect 450 128 451 132
rect 411 84 451 128
rect 455 4055 461 4172
rect 455 4051 456 4055
rect 460 4051 461 4055
rect 455 4045 461 4051
rect 455 4041 456 4045
rect 460 4041 461 4045
rect 455 4017 461 4041
rect 455 4013 456 4017
rect 460 4013 461 4017
rect 455 4007 461 4013
rect 455 4003 456 4007
rect 460 4003 461 4007
rect 455 3581 461 4003
rect 455 3577 456 3581
rect 460 3577 461 3581
rect 455 3571 461 3577
rect 455 3567 456 3571
rect 460 3567 461 3571
rect 455 3543 461 3567
rect 455 3539 456 3543
rect 460 3539 461 3543
rect 455 3533 461 3539
rect 455 3529 456 3533
rect 460 3529 461 3533
rect 455 3107 461 3529
rect 455 3103 456 3107
rect 460 3103 461 3107
rect 455 3097 461 3103
rect 455 3093 456 3097
rect 460 3093 461 3097
rect 455 3069 461 3093
rect 455 3065 456 3069
rect 460 3065 461 3069
rect 455 3059 461 3065
rect 455 3055 456 3059
rect 460 3055 461 3059
rect 455 2633 461 3055
rect 455 2629 456 2633
rect 460 2629 461 2633
rect 455 2623 461 2629
rect 455 2619 456 2623
rect 460 2619 461 2623
rect 455 2595 461 2619
rect 455 2591 456 2595
rect 460 2591 461 2595
rect 455 2585 461 2591
rect 455 2581 456 2585
rect 460 2581 461 2585
rect 455 2159 461 2581
rect 455 2155 456 2159
rect 460 2155 461 2159
rect 455 2149 461 2155
rect 455 2145 456 2149
rect 460 2145 461 2149
rect 455 2121 461 2145
rect 455 2117 456 2121
rect 460 2117 461 2121
rect 455 2111 461 2117
rect 455 2107 456 2111
rect 460 2107 461 2111
rect 455 1685 461 2107
rect 455 1681 456 1685
rect 460 1681 461 1685
rect 455 1675 461 1681
rect 455 1671 456 1675
rect 460 1671 461 1675
rect 455 1647 461 1671
rect 455 1643 456 1647
rect 460 1643 461 1647
rect 455 1637 461 1643
rect 455 1633 456 1637
rect 460 1633 461 1637
rect 455 1211 461 1633
rect 455 1207 456 1211
rect 460 1207 461 1211
rect 455 1201 461 1207
rect 455 1197 456 1201
rect 460 1197 461 1201
rect 455 1173 461 1197
rect 455 1169 456 1173
rect 460 1169 461 1173
rect 455 1163 461 1169
rect 455 1159 456 1163
rect 460 1159 461 1163
rect 455 737 461 1159
rect 455 733 456 737
rect 460 733 461 737
rect 455 727 461 733
rect 455 723 456 727
rect 460 723 461 727
rect 455 699 461 723
rect 455 695 456 699
rect 460 695 461 699
rect 455 689 461 695
rect 455 685 456 689
rect 460 685 461 689
rect 455 263 461 685
rect 455 259 456 263
rect 460 259 461 263
rect 455 253 461 259
rect 455 249 456 253
rect 460 249 461 253
rect 455 225 461 249
rect 455 221 456 225
rect 460 221 461 225
rect 455 215 461 221
rect 455 211 456 215
rect 460 211 461 215
rect 455 94 461 211
rect 465 4094 505 4168
rect 465 4090 466 4094
rect 470 4090 477 4094
rect 481 4090 483 4094
rect 487 4090 495 4094
rect 499 4090 509 4094
rect 465 4088 513 4090
rect 465 4084 466 4088
rect 470 4084 477 4088
rect 481 4084 483 4088
rect 487 4084 495 4088
rect 499 4084 509 4088
rect 465 4082 513 4084
rect 465 4078 466 4082
rect 470 4078 477 4082
rect 481 4078 483 4082
rect 487 4078 495 4082
rect 499 4078 509 4082
rect 465 4076 513 4078
rect 465 4072 466 4076
rect 470 4072 477 4076
rect 481 4072 483 4076
rect 487 4072 495 4076
rect 499 4072 509 4076
rect 465 4070 513 4072
rect 465 4066 466 4070
rect 470 4066 477 4070
rect 481 4066 483 4070
rect 487 4066 495 4070
rect 499 4066 509 4070
rect 465 4064 513 4066
rect 465 4060 466 4064
rect 470 4060 477 4064
rect 481 4060 483 4064
rect 487 4060 495 4064
rect 499 4060 509 4064
rect 465 4058 513 4060
rect 465 4054 466 4058
rect 470 4054 477 4058
rect 481 4054 483 4058
rect 487 4054 495 4058
rect 499 4054 509 4058
rect 465 4004 505 4054
rect 465 4000 466 4004
rect 470 4000 477 4004
rect 481 4000 483 4004
rect 487 4000 495 4004
rect 499 4000 509 4004
rect 465 3998 513 4000
rect 465 3994 466 3998
rect 470 3994 477 3998
rect 481 3994 483 3998
rect 487 3994 495 3998
rect 499 3994 509 3998
rect 465 3992 513 3994
rect 465 3988 466 3992
rect 470 3988 477 3992
rect 481 3988 483 3992
rect 487 3988 495 3992
rect 499 3988 509 3992
rect 465 3986 513 3988
rect 465 3982 466 3986
rect 470 3982 477 3986
rect 481 3982 483 3986
rect 487 3982 495 3986
rect 499 3982 509 3986
rect 465 3980 513 3982
rect 465 3976 466 3980
rect 470 3976 477 3980
rect 481 3976 483 3980
rect 487 3976 495 3980
rect 499 3976 509 3980
rect 465 3974 513 3976
rect 465 3970 466 3974
rect 470 3970 477 3974
rect 481 3970 483 3974
rect 487 3970 495 3974
rect 499 3970 509 3974
rect 465 3968 513 3970
rect 465 3964 466 3968
rect 470 3964 477 3968
rect 481 3964 483 3968
rect 487 3964 509 3968
rect 465 3620 505 3964
rect 509 3954 513 3956
rect 509 3948 513 3950
rect 509 3942 513 3944
rect 509 3936 513 3938
rect 509 3930 513 3932
rect 509 3924 513 3926
rect 509 3658 513 3660
rect 509 3652 513 3654
rect 509 3646 513 3648
rect 509 3640 513 3642
rect 509 3634 513 3636
rect 509 3628 513 3630
rect 469 3616 477 3620
rect 481 3616 483 3620
rect 487 3616 509 3620
rect 465 3614 513 3616
rect 469 3610 477 3614
rect 481 3610 483 3614
rect 487 3610 495 3614
rect 499 3610 509 3614
rect 465 3608 513 3610
rect 469 3604 477 3608
rect 481 3604 483 3608
rect 487 3604 495 3608
rect 499 3604 509 3608
rect 465 3602 513 3604
rect 469 3598 477 3602
rect 481 3598 483 3602
rect 487 3598 495 3602
rect 499 3598 509 3602
rect 465 3596 513 3598
rect 469 3592 477 3596
rect 481 3592 483 3596
rect 487 3592 495 3596
rect 499 3592 509 3596
rect 465 3590 513 3592
rect 469 3586 477 3590
rect 481 3586 483 3590
rect 487 3586 495 3590
rect 499 3586 509 3590
rect 465 3584 513 3586
rect 469 3580 477 3584
rect 481 3580 483 3584
rect 487 3580 495 3584
rect 499 3580 509 3584
rect 465 3530 505 3580
rect 469 3526 477 3530
rect 481 3526 483 3530
rect 487 3526 495 3530
rect 499 3526 509 3530
rect 465 3524 513 3526
rect 469 3520 477 3524
rect 481 3520 483 3524
rect 487 3520 495 3524
rect 499 3520 509 3524
rect 465 3518 513 3520
rect 469 3514 477 3518
rect 481 3514 483 3518
rect 487 3514 495 3518
rect 499 3514 509 3518
rect 465 3512 513 3514
rect 469 3508 477 3512
rect 481 3508 483 3512
rect 487 3508 495 3512
rect 499 3508 509 3512
rect 465 3506 513 3508
rect 469 3502 477 3506
rect 481 3502 483 3506
rect 487 3502 495 3506
rect 499 3502 509 3506
rect 465 3500 513 3502
rect 469 3496 477 3500
rect 481 3496 483 3500
rect 487 3496 495 3500
rect 499 3496 509 3500
rect 465 3494 513 3496
rect 469 3490 477 3494
rect 481 3490 483 3494
rect 487 3490 509 3494
rect 465 3146 505 3490
rect 509 3480 513 3482
rect 509 3474 513 3476
rect 509 3468 513 3470
rect 509 3462 513 3464
rect 509 3456 513 3458
rect 509 3450 513 3452
rect 509 3184 513 3186
rect 509 3178 513 3180
rect 509 3172 513 3174
rect 509 3166 513 3168
rect 509 3160 513 3162
rect 509 3154 513 3156
rect 469 3142 477 3146
rect 481 3142 483 3146
rect 487 3142 509 3146
rect 465 3140 513 3142
rect 469 3136 477 3140
rect 481 3136 483 3140
rect 487 3136 495 3140
rect 499 3136 509 3140
rect 465 3134 513 3136
rect 469 3130 477 3134
rect 481 3130 483 3134
rect 487 3130 495 3134
rect 499 3130 509 3134
rect 465 3128 513 3130
rect 469 3124 477 3128
rect 481 3124 483 3128
rect 487 3124 495 3128
rect 499 3124 509 3128
rect 465 3122 513 3124
rect 469 3118 477 3122
rect 481 3118 483 3122
rect 487 3118 495 3122
rect 499 3118 509 3122
rect 465 3116 513 3118
rect 469 3112 477 3116
rect 481 3112 483 3116
rect 487 3112 495 3116
rect 499 3112 509 3116
rect 465 3110 513 3112
rect 469 3106 477 3110
rect 481 3106 483 3110
rect 487 3106 495 3110
rect 499 3106 509 3110
rect 465 3056 505 3106
rect 469 3052 477 3056
rect 481 3052 483 3056
rect 487 3052 495 3056
rect 499 3052 509 3056
rect 465 3050 513 3052
rect 469 3046 477 3050
rect 481 3046 483 3050
rect 487 3046 495 3050
rect 499 3046 509 3050
rect 465 3044 513 3046
rect 469 3040 477 3044
rect 481 3040 483 3044
rect 487 3040 495 3044
rect 499 3040 509 3044
rect 465 3038 513 3040
rect 469 3034 477 3038
rect 481 3034 483 3038
rect 487 3034 495 3038
rect 499 3034 509 3038
rect 465 3032 513 3034
rect 469 3028 477 3032
rect 481 3028 483 3032
rect 487 3028 495 3032
rect 499 3028 509 3032
rect 465 3026 513 3028
rect 469 3022 477 3026
rect 481 3022 483 3026
rect 487 3022 495 3026
rect 499 3022 509 3026
rect 465 3020 513 3022
rect 469 3016 477 3020
rect 481 3016 483 3020
rect 487 3016 509 3020
rect 465 2672 505 3016
rect 509 3006 513 3008
rect 509 3000 513 3002
rect 509 2994 513 2996
rect 509 2988 513 2990
rect 509 2982 513 2984
rect 509 2976 513 2978
rect 509 2710 513 2712
rect 509 2704 513 2706
rect 509 2698 513 2700
rect 509 2692 513 2694
rect 509 2686 513 2688
rect 509 2680 513 2682
rect 469 2668 477 2672
rect 481 2668 483 2672
rect 487 2668 509 2672
rect 465 2666 513 2668
rect 469 2662 477 2666
rect 481 2662 483 2666
rect 487 2662 495 2666
rect 499 2662 509 2666
rect 465 2660 513 2662
rect 469 2656 477 2660
rect 481 2656 483 2660
rect 487 2656 495 2660
rect 499 2656 509 2660
rect 465 2654 513 2656
rect 469 2650 477 2654
rect 481 2650 483 2654
rect 487 2650 495 2654
rect 499 2650 509 2654
rect 465 2648 513 2650
rect 469 2644 477 2648
rect 481 2644 483 2648
rect 487 2644 495 2648
rect 499 2644 509 2648
rect 465 2642 513 2644
rect 469 2638 477 2642
rect 481 2638 483 2642
rect 487 2638 495 2642
rect 499 2638 509 2642
rect 465 2636 513 2638
rect 469 2632 477 2636
rect 481 2632 483 2636
rect 487 2632 495 2636
rect 499 2632 509 2636
rect 465 2582 505 2632
rect 469 2578 477 2582
rect 481 2578 483 2582
rect 487 2578 495 2582
rect 499 2578 509 2582
rect 465 2576 513 2578
rect 469 2572 477 2576
rect 481 2572 483 2576
rect 487 2572 495 2576
rect 499 2572 509 2576
rect 465 2570 513 2572
rect 469 2566 477 2570
rect 481 2566 483 2570
rect 487 2566 495 2570
rect 499 2566 509 2570
rect 465 2564 513 2566
rect 469 2560 477 2564
rect 481 2560 483 2564
rect 487 2560 495 2564
rect 499 2560 509 2564
rect 465 2558 513 2560
rect 469 2554 477 2558
rect 481 2554 483 2558
rect 487 2554 495 2558
rect 499 2554 509 2558
rect 465 2552 513 2554
rect 469 2548 477 2552
rect 481 2548 483 2552
rect 487 2548 495 2552
rect 499 2548 509 2552
rect 465 2546 513 2548
rect 469 2542 477 2546
rect 481 2542 483 2546
rect 487 2542 509 2546
rect 465 2198 505 2542
rect 509 2532 513 2534
rect 509 2526 513 2528
rect 509 2520 513 2522
rect 509 2514 513 2516
rect 509 2508 513 2510
rect 509 2502 513 2504
rect 509 2236 513 2238
rect 509 2230 513 2232
rect 509 2224 513 2226
rect 509 2218 513 2220
rect 509 2212 513 2214
rect 509 2206 513 2208
rect 469 2194 477 2198
rect 481 2194 483 2198
rect 487 2194 509 2198
rect 465 2192 513 2194
rect 469 2188 477 2192
rect 481 2188 483 2192
rect 487 2188 495 2192
rect 499 2188 509 2192
rect 465 2186 513 2188
rect 469 2182 477 2186
rect 481 2182 483 2186
rect 487 2182 495 2186
rect 499 2182 509 2186
rect 465 2180 513 2182
rect 469 2176 477 2180
rect 481 2176 483 2180
rect 487 2176 495 2180
rect 499 2176 509 2180
rect 465 2174 513 2176
rect 469 2170 477 2174
rect 481 2170 483 2174
rect 487 2170 495 2174
rect 499 2170 509 2174
rect 465 2168 513 2170
rect 469 2164 477 2168
rect 481 2164 483 2168
rect 487 2164 495 2168
rect 499 2164 509 2168
rect 465 2162 513 2164
rect 469 2158 477 2162
rect 481 2158 483 2162
rect 487 2158 495 2162
rect 499 2158 509 2162
rect 465 2108 505 2158
rect 469 2104 477 2108
rect 481 2104 483 2108
rect 487 2104 495 2108
rect 499 2104 509 2108
rect 465 2102 513 2104
rect 469 2098 477 2102
rect 481 2098 483 2102
rect 487 2098 495 2102
rect 499 2098 509 2102
rect 465 2096 513 2098
rect 469 2092 477 2096
rect 481 2092 483 2096
rect 487 2092 495 2096
rect 499 2092 509 2096
rect 465 2090 513 2092
rect 469 2086 477 2090
rect 481 2086 483 2090
rect 487 2086 495 2090
rect 499 2086 509 2090
rect 465 2084 513 2086
rect 469 2080 477 2084
rect 481 2080 483 2084
rect 487 2080 495 2084
rect 499 2080 509 2084
rect 465 2078 513 2080
rect 469 2074 477 2078
rect 481 2074 483 2078
rect 487 2074 495 2078
rect 499 2074 509 2078
rect 465 2072 513 2074
rect 469 2068 477 2072
rect 481 2068 483 2072
rect 487 2068 509 2072
rect 465 1724 505 2068
rect 509 2058 513 2060
rect 509 2052 513 2054
rect 509 2046 513 2048
rect 509 2040 513 2042
rect 509 2034 513 2036
rect 509 2028 513 2030
rect 509 1762 513 1764
rect 509 1756 513 1758
rect 509 1750 513 1752
rect 509 1744 513 1746
rect 509 1738 513 1740
rect 509 1732 513 1734
rect 469 1720 477 1724
rect 481 1720 483 1724
rect 487 1720 509 1724
rect 465 1718 513 1720
rect 469 1714 477 1718
rect 481 1714 483 1718
rect 487 1714 495 1718
rect 499 1714 509 1718
rect 465 1712 513 1714
rect 469 1708 477 1712
rect 481 1708 483 1712
rect 487 1708 495 1712
rect 499 1708 509 1712
rect 465 1706 513 1708
rect 469 1702 477 1706
rect 481 1702 483 1706
rect 487 1702 495 1706
rect 499 1702 509 1706
rect 465 1700 513 1702
rect 469 1696 477 1700
rect 481 1696 483 1700
rect 487 1696 495 1700
rect 499 1696 509 1700
rect 465 1694 513 1696
rect 469 1690 477 1694
rect 481 1690 483 1694
rect 487 1690 495 1694
rect 499 1690 509 1694
rect 465 1688 513 1690
rect 469 1684 477 1688
rect 481 1684 483 1688
rect 487 1684 495 1688
rect 499 1684 509 1688
rect 465 1634 505 1684
rect 469 1630 477 1634
rect 481 1630 483 1634
rect 487 1630 495 1634
rect 499 1630 509 1634
rect 465 1628 513 1630
rect 469 1624 477 1628
rect 481 1624 483 1628
rect 487 1624 495 1628
rect 499 1624 509 1628
rect 465 1622 513 1624
rect 469 1618 477 1622
rect 481 1618 483 1622
rect 487 1618 495 1622
rect 499 1618 509 1622
rect 465 1616 513 1618
rect 469 1612 477 1616
rect 481 1612 483 1616
rect 487 1612 495 1616
rect 499 1612 509 1616
rect 465 1610 513 1612
rect 469 1606 477 1610
rect 481 1606 483 1610
rect 487 1606 495 1610
rect 499 1606 509 1610
rect 465 1604 513 1606
rect 469 1600 477 1604
rect 481 1600 483 1604
rect 487 1600 495 1604
rect 499 1600 509 1604
rect 465 1598 513 1600
rect 469 1594 477 1598
rect 481 1594 483 1598
rect 487 1594 509 1598
rect 465 1250 505 1594
rect 509 1584 513 1586
rect 509 1578 513 1580
rect 509 1572 513 1574
rect 509 1566 513 1568
rect 509 1560 513 1562
rect 509 1554 513 1556
rect 509 1288 513 1290
rect 509 1282 513 1284
rect 509 1276 513 1278
rect 509 1270 513 1272
rect 509 1264 513 1266
rect 509 1258 513 1260
rect 469 1246 477 1250
rect 481 1246 483 1250
rect 487 1246 509 1250
rect 465 1244 513 1246
rect 469 1240 477 1244
rect 481 1240 483 1244
rect 487 1240 495 1244
rect 499 1240 509 1244
rect 465 1238 513 1240
rect 469 1234 477 1238
rect 481 1234 483 1238
rect 487 1234 495 1238
rect 499 1234 509 1238
rect 465 1232 513 1234
rect 469 1228 477 1232
rect 481 1228 483 1232
rect 487 1228 495 1232
rect 499 1228 509 1232
rect 465 1226 513 1228
rect 469 1222 477 1226
rect 481 1222 483 1226
rect 487 1222 495 1226
rect 499 1222 509 1226
rect 465 1220 513 1222
rect 469 1216 477 1220
rect 481 1216 483 1220
rect 487 1216 495 1220
rect 499 1216 509 1220
rect 465 1214 513 1216
rect 469 1210 477 1214
rect 481 1210 483 1214
rect 487 1210 495 1214
rect 499 1210 509 1214
rect 465 1160 505 1210
rect 469 1156 477 1160
rect 481 1156 483 1160
rect 487 1156 495 1160
rect 499 1156 509 1160
rect 465 1154 513 1156
rect 469 1150 477 1154
rect 481 1150 483 1154
rect 487 1150 495 1154
rect 499 1150 509 1154
rect 465 1148 513 1150
rect 469 1144 477 1148
rect 481 1144 483 1148
rect 487 1144 495 1148
rect 499 1144 509 1148
rect 465 1142 513 1144
rect 469 1138 477 1142
rect 481 1138 483 1142
rect 487 1138 495 1142
rect 499 1138 509 1142
rect 465 1136 513 1138
rect 469 1132 477 1136
rect 481 1132 483 1136
rect 487 1132 495 1136
rect 499 1132 509 1136
rect 465 1130 513 1132
rect 469 1126 477 1130
rect 481 1126 483 1130
rect 487 1126 495 1130
rect 499 1126 509 1130
rect 465 1124 513 1126
rect 469 1120 477 1124
rect 481 1120 483 1124
rect 487 1120 509 1124
rect 465 776 505 1120
rect 509 1110 513 1112
rect 509 1104 513 1106
rect 509 1098 513 1100
rect 509 1092 513 1094
rect 509 1086 513 1088
rect 509 1080 513 1082
rect 509 814 513 816
rect 509 808 513 810
rect 509 802 513 804
rect 509 796 513 798
rect 509 790 513 792
rect 509 784 513 786
rect 469 772 477 776
rect 481 772 483 776
rect 487 772 509 776
rect 465 770 513 772
rect 469 766 477 770
rect 481 766 483 770
rect 487 766 495 770
rect 499 766 509 770
rect 465 764 513 766
rect 469 760 477 764
rect 481 760 483 764
rect 487 760 495 764
rect 499 760 509 764
rect 465 758 513 760
rect 469 754 477 758
rect 481 754 483 758
rect 487 754 495 758
rect 499 754 509 758
rect 465 752 513 754
rect 469 748 477 752
rect 481 748 483 752
rect 487 748 495 752
rect 499 748 509 752
rect 465 746 513 748
rect 469 742 477 746
rect 481 742 483 746
rect 487 742 495 746
rect 499 742 509 746
rect 465 740 513 742
rect 469 736 477 740
rect 481 736 483 740
rect 487 736 495 740
rect 499 736 509 740
rect 465 686 505 736
rect 469 682 477 686
rect 481 682 483 686
rect 487 682 495 686
rect 499 682 509 686
rect 465 680 513 682
rect 469 676 477 680
rect 481 676 483 680
rect 487 676 495 680
rect 499 676 509 680
rect 465 674 513 676
rect 469 670 477 674
rect 481 670 483 674
rect 487 670 495 674
rect 499 670 509 674
rect 465 668 513 670
rect 469 664 477 668
rect 481 664 483 668
rect 487 664 495 668
rect 499 664 509 668
rect 465 662 513 664
rect 469 658 477 662
rect 481 658 483 662
rect 487 658 495 662
rect 499 658 509 662
rect 465 656 513 658
rect 469 652 477 656
rect 481 652 483 656
rect 487 652 495 656
rect 499 652 509 656
rect 465 650 513 652
rect 469 646 477 650
rect 481 646 483 650
rect 487 646 509 650
rect 465 302 505 646
rect 509 636 513 638
rect 509 630 513 632
rect 509 624 513 626
rect 509 618 513 620
rect 509 612 513 614
rect 509 606 513 608
rect 509 340 513 342
rect 509 334 513 336
rect 509 328 513 330
rect 509 322 513 324
rect 509 316 513 318
rect 509 310 513 312
rect 469 298 477 302
rect 481 298 483 302
rect 487 298 509 302
rect 465 296 513 298
rect 469 292 477 296
rect 481 292 483 296
rect 487 292 495 296
rect 499 292 509 296
rect 465 290 513 292
rect 469 286 477 290
rect 481 286 483 290
rect 487 286 495 290
rect 499 286 509 290
rect 465 284 513 286
rect 469 280 477 284
rect 481 280 483 284
rect 487 280 495 284
rect 499 280 509 284
rect 465 278 513 280
rect 469 274 477 278
rect 481 274 483 278
rect 487 274 495 278
rect 499 274 509 278
rect 465 272 513 274
rect 469 268 477 272
rect 481 268 483 272
rect 487 268 495 272
rect 499 268 509 272
rect 465 266 513 268
rect 469 262 477 266
rect 481 262 483 266
rect 487 262 495 266
rect 499 262 509 266
rect 465 212 505 262
rect 469 208 477 212
rect 481 208 483 212
rect 487 208 495 212
rect 499 208 509 212
rect 465 206 513 208
rect 469 202 477 206
rect 481 202 483 206
rect 487 202 495 206
rect 499 202 509 206
rect 465 200 513 202
rect 469 196 477 200
rect 481 196 483 200
rect 487 196 495 200
rect 499 196 509 200
rect 465 194 513 196
rect 469 190 477 194
rect 481 190 483 194
rect 487 190 495 194
rect 499 190 509 194
rect 465 188 513 190
rect 469 184 477 188
rect 481 184 483 188
rect 487 184 495 188
rect 499 184 509 188
rect 465 182 513 184
rect 469 178 477 182
rect 481 178 483 182
rect 487 178 495 182
rect 499 178 509 182
rect 465 176 513 178
rect 469 172 477 176
rect 481 172 483 176
rect 487 172 495 176
rect 499 172 509 176
rect 465 164 505 172
rect 465 135 467 164
rect 496 135 505 164
rect 465 98 505 135
<< m3contact >>
rect 413 4146 447 4180
rect 467 135 496 164
<< metal3 >>
rect 412 4180 448 4184
rect 412 4146 413 4180
rect 447 4146 448 4180
rect 412 4145 448 4146
rect 466 164 497 165
rect 466 135 467 164
rect 496 135 497 164
rect 466 130 497 135
<< labels >>
rlabel m2contact 512 326 512 326 6 Gnd
rlabel m2contact 512 192 512 192 6 CVdd
rlabel m2contact 512 220 512 220 6 Bias
rlabel m2contact 512 253 512 253 6 Bias
rlabel m2contact 512 282 512 282 6 CVdd
rlabel m2contact 512 800 512 800 6 Gnd
rlabel m2contact 512 622 512 622 6 Gnd
rlabel m2contact 512 666 512 666 6 CVdd
rlabel m2contact 512 694 512 694 6 Bias
rlabel m2contact 512 727 512 727 6 Bias
rlabel m2contact 512 756 512 756 6 CVdd
rlabel m2contact 512 1274 512 1274 6 Gnd
rlabel m2contact 512 1096 512 1096 6 Gnd
rlabel m2contact 512 1140 512 1140 6 CVdd
rlabel m2contact 512 1168 512 1168 6 Bias
rlabel m2contact 512 1201 512 1201 6 Bias
rlabel m2contact 512 1230 512 1230 6 CVdd
rlabel m2contact 512 1748 512 1748 6 Gnd
rlabel m2contact 512 1570 512 1570 6 Gnd
rlabel m2contact 512 1614 512 1614 6 CVdd
rlabel m2contact 512 1642 512 1642 6 Bias
rlabel m2contact 512 1675 512 1675 6 Bias
rlabel m2contact 512 1704 512 1704 6 CVdd
rlabel m2contact 512 2222 512 2222 6 Gnd
rlabel m2contact 512 2044 512 2044 6 Gnd
rlabel m2contact 512 2088 512 2088 6 CVdd
rlabel m2contact 512 2116 512 2116 6 Bias
rlabel m2contact 512 2149 512 2149 6 Bias
rlabel m2contact 512 2178 512 2178 6 CVdd
rlabel m2contact 512 2696 512 2696 6 Gnd
rlabel m2contact 512 2518 512 2518 6 Gnd
rlabel m2contact 512 2562 512 2562 6 CVdd
rlabel m2contact 512 2590 512 2590 6 Bias
rlabel m2contact 512 2623 512 2623 6 Bias
rlabel m2contact 512 2652 512 2652 6 CVdd
rlabel m2contact 512 3170 512 3170 6 Gnd
rlabel m2contact 512 2992 512 2992 6 Gnd
rlabel m2contact 512 3036 512 3036 6 CVdd
rlabel m2contact 512 3064 512 3064 6 Bias
rlabel m2contact 512 3097 512 3097 6 Bias
rlabel m2contact 512 3126 512 3126 6 CVdd
rlabel m2contact 512 3644 512 3644 6 Gnd
rlabel m2contact 512 3466 512 3466 6 Gnd
rlabel m2contact 512 3510 512 3510 6 CVdd
rlabel m2contact 512 3538 512 3538 6 Bias
rlabel m2contact 512 3571 512 3571 6 Bias
rlabel m2contact 512 3600 512 3600 6 CVdd
rlabel m2contact 512 3940 512 3940 6 Gnd
rlabel m2contact 512 3984 512 3984 6 CVdd
rlabel m2contact 512 4012 512 4012 6 Bias
rlabel m2contact 512 4045 512 4045 6 Bias
rlabel m2contact 512 4074 512 4074 6 CVdd
<< end >>
