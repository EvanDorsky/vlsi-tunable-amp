magic
tech scmos
timestamp 1418704018
<< ntransistor >>
rect 0 0 6 120
rect 0 -129 6 -9
<< ptransistor >>
rect -24 0 -18 120
rect -24 -129 -18 -9
<< ndiffusion >>
rect -3 0 0 120
rect 6 4 9 120
rect 6 0 7 4
rect -3 -129 0 -9
rect 6 -13 7 -9
rect 6 -129 9 -13
<< pdiffusion >>
rect -27 4 -24 120
rect -25 0 -24 4
rect -18 0 -15 120
rect -25 -13 -24 -9
rect -27 -129 -24 -13
rect -18 -129 -15 -9
<< ndcontact >>
rect 7 0 11 4
rect 7 -13 11 -9
<< pdcontact >>
rect -29 0 -25 4
rect -29 -13 -25 -9
<< polysilicon >>
rect -24 120 -18 123
rect 0 120 6 123
rect -24 -1 -18 0
rect 0 -1 6 0
rect -24 -3 6 -1
rect -24 -8 6 -6
rect -24 -9 -18 -8
rect 0 -9 6 -8
rect -24 -132 -18 -129
rect 0 -132 6 -129
<< metal1 >>
rect -29 -9 -25 0
rect 7 -9 11 0
<< labels >>
rlabel metal1 7 -9 11 0 3 Gnd
rlabel metal1 -29 -9 -25 0 3 Vdd
rlabel polysilicon -18 -8 0 -6 1 V-
rlabel polysilicon -18 -3 0 -1 1 V+
<< end >>
