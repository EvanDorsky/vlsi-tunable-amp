magic
tech scmos
timestamp 1418873168
use barepad  barepad_1
timestamp 1259953556
transform -1 0 841 0 -1 5000
box -2 0 476 513
use inpad  inpad_1
timestamp 1259953556
transform -1 0 1315 0 -1 5000
box -2 0 476 513
use inpad  inpad_0
timestamp 1259953556
transform -1 0 1789 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_3
timestamp 1259953556
transform -1 0 2263 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_6
timestamp 1259953556
transform -1 0 2737 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_5
timestamp 1259953556
transform -1 0 3211 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_4
timestamp 1259953556
transform -1 0 3685 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_3
timestamp 1259953556
transform -1 0 4159 0 -1 5000
box -2 0 476 513
use barepad  barepad_0
timestamp 1259953556
transform -1 0 4633 0 -1 5000
box -2 0 476 513
use padframe_top  padframe_top_0
timestamp 1259953556
transform 1 0 0 0 1 4487
box 0 0 5000 513
use barepad  barepad_2
timestamp 1259953556
transform 0 1 0 -1 0 4633
box -2 0 476 513
use inorpad  inorpad_7
timestamp 1259953556
transform 0 1 0 -1 0 4159
box -2 0 476 513
use inorpad  inorpad_8
timestamp 1259953556
transform 0 1 0 -1 0 3685
box -2 0 476 513
use inorpad  inorpad_9
timestamp 1259953556
transform 0 1 0 -1 0 3211
box -2 0 476 513
use inorpad  inorpad_10
timestamp 1259953556
transform 0 1 0 -1 0 2737
box -2 0 476 513
use inpad  inpad_2
timestamp 1259953556
transform 0 1 0 -1 0 2263
box -2 0 476 513
use inpad  inpad_3
timestamp 1259953556
transform 0 1 0 -1 0 1789
box -2 0 476 513
use inpad  inpad_4
timestamp 1259953556
transform 0 1 0 -1 0 1315
box -2 0 476 513
use inorpad  inorpad_17
timestamp 1259953556
transform 0 -1 5000 1 0 4159
box -2 0 476 513
use inorpad  inorpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 3685
box -2 0 476 513
use inorpad  inorpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 3211
box -2 0 476 513
use inorpad  inorpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 2737
box -2 0 476 513
use blankpad  blankpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 2263
box -2 0 476 513
use blankpad  blankpad_7
timestamp 1259953556
transform 0 -1 5000 1 0 1789
box -2 0 476 513
use blankpad  blankpad_8
timestamp 1259953556
transform 0 -1 5000 1 0 1315
box -2 0 476 513
use blankpad  blankpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 841
box -2 0 476 513
use padframe_left  padframe_left_0
timestamp 1259953556
transform 1 0 0 0 1 367
box 2 2 513 4264
use iopad  iopad_0
timestamp 1259953556
transform 0 1 0 -1 0 841
box -2 0 476 513
use iopad  iopad_1
timestamp 1259953556
transform 1 0 367 0 1 0
box -2 0 476 513
use inorpad  inorpad_11
timestamp 1259953556
transform 1 0 841 0 1 0
box -2 0 476 513
use inorpad  inorpad_12
timestamp 1259953556
transform 1 0 1315 0 1 0
box -2 0 476 513
use iopad  iopad_2
timestamp 1259953556
transform 1 0 1789 0 1 0
box -2 0 476 513
use iopad  iopad_3
timestamp 1259953556
transform 1 0 2263 0 1 0
box -2 0 476 513
use inorpad  inorpad_13
timestamp 1259953556
transform 1 0 2737 0 1 0
box -2 0 476 513
use inorpad  inorpad_14
timestamp 1259953556
transform 1 0 3211 0 1 0
box -2 0 476 513
use inorpad  inorpad_15
timestamp 1259953556
transform 1 0 3685 0 1 0
box -2 0 476 513
use padframe_right  padframe_right_0
timestamp 1259953556
transform 1 0 4487 0 1 367
box 0 2 511 4264
use blankpad  blankpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 367
box -2 0 476 513
use inorpad  inorpad_16
timestamp 1259953556
transform 1 0 4159 0 1 0
box -2 0 476 513
use padframe_bottom  padframe_bottom_0
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 5000 513
<< end >>
