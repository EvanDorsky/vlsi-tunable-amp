magic
tech scmos
magscale 1 3
timestamp 1419146600
<< nwell >>
rect 4668 4263 4680 4275
rect 4971 4203 5028 4281
rect 2571 3600 2622 3849
rect 8241 3846 8316 3849
rect 8241 3840 8325 3846
rect 8241 3600 8292 3840
rect 8274 3597 8292 3600
<< nsubstratencontact >>
rect 2586 3696 2607 3828
rect 8256 3696 8277 3828
<< polysilicon >>
rect 4017 4302 5028 4335
rect 4017 4206 4056 4302
rect 4668 4263 4680 4272
rect 4989 4251 5028 4302
rect 10335 4260 10347 4269
rect 7020 3087 7032 3099
rect 12720 3087 12732 3099
<< polycontact >>
rect 3588 4206 3600 4218
rect 4668 4272 4680 4284
rect 10335 4269 10347 4281
rect 4989 4203 5028 4251
rect 9258 4203 9276 4215
rect 7008 3087 7020 3099
rect 7032 3087 7044 3099
rect 12708 3087 12720 3099
rect 12732 3087 12744 3099
<< metal1 >>
rect 2214 4413 2274 4422
rect 7881 4410 7890 4587
rect 4524 4317 4578 4320
rect 4323 4311 4578 4317
rect 4323 4308 4548 4311
rect 4590 4311 4599 4320
rect 10095 4317 10107 4344
rect 3666 4302 3924 4305
rect 4323 4302 4335 4308
rect 10269 4317 10281 4347
rect 3666 4299 4335 4302
rect 3429 4293 4335 4299
rect 3429 4287 3675 4293
rect 7116 4266 7140 4275
rect 3327 4161 3348 4245
rect 3462 4242 3468 4254
rect 3492 4242 3498 4254
rect 5118 4260 7140 4266
rect 5118 4254 7125 4260
rect 7173 4254 7182 4281
rect 7218 4257 7251 4275
rect 3462 4104 3498 4242
rect 5073 4230 7140 4242
rect 7173 4230 7182 4251
rect 7239 4248 9285 4257
rect 7218 4239 7230 4242
rect 7218 4236 9276 4239
rect 7218 4230 9318 4236
rect 7227 4227 9318 4230
rect 5028 4203 7140 4221
rect 7218 4203 9258 4215
rect 3495 4077 3498 4104
rect 3462 4074 3498 4077
rect 7638 3894 7743 3897
rect 1665 3849 2607 3894
rect 7638 3849 8277 3894
rect 1665 3840 2673 3849
rect 7638 3846 8316 3849
rect 7638 3840 8358 3846
rect 1665 3834 2607 3840
rect 1665 2010 1737 3834
rect 2586 3828 2607 3834
rect 7638 3834 8277 3840
rect 8307 3837 8358 3840
rect 7638 3306 7743 3834
rect 8256 3828 8277 3834
rect 6777 3081 6951 3111
rect 6777 3066 6858 3081
rect 7008 3075 7044 3087
rect 7635 2820 7743 3306
rect 12423 3099 12522 3108
rect 12423 3087 12432 3099
rect 12444 3063 12522 3099
rect 12708 3075 12744 3087
rect 2208 2304 2637 2328
rect 1527 1887 1737 2010
rect 1665 1869 1737 1887
rect 1554 1833 1737 1869
rect 1527 1791 1737 1833
rect 1554 1761 1737 1791
rect 1668 1737 1737 1761
rect 1527 1614 1737 1737
rect 1788 2283 3948 2286
rect 7635 2283 7740 2820
rect 1788 2229 7740 2283
rect 1788 2193 7734 2229
rect 1788 1614 1833 2193
rect 3837 2190 7734 2193
rect 1788 1599 2007 1614
rect 1617 1572 2007 1599
rect 1617 1566 1833 1572
rect 1617 1527 1737 1566
rect 1788 1527 1833 1566
rect 1887 1527 2007 1572
<< m2contact >>
rect 7881 4587 7893 4599
rect 2274 4413 2286 4425
rect 10095 4344 10107 4356
rect 4578 4308 4590 4320
rect 10095 4305 10107 4317
rect 10269 4347 10281 4359
rect 10269 4305 10281 4317
rect 3417 4287 3429 4299
rect 4656 4272 4668 4284
rect 3327 4245 3357 4260
rect 3468 4242 3492 4260
rect 3780 4251 3792 4263
rect 3852 4251 3864 4263
rect 5103 4254 5118 4266
rect 7140 4257 7158 4275
rect 7200 4257 7218 4275
rect 10323 4269 10335 4281
rect 3324 4134 3357 4161
rect 3576 4206 3588 4218
rect 5058 4230 5073 4242
rect 7140 4230 7158 4248
rect 7200 4230 7218 4248
rect 9285 4245 9300 4257
rect 9318 4227 9333 4242
rect 7140 4203 7158 4221
rect 7200 4203 7218 4221
rect 3462 4077 3495 4104
rect 6858 3051 6951 3081
rect 7008 3063 7044 3075
rect 12522 3063 12621 3108
rect 12708 3063 12744 3075
rect 2148 2304 2208 2328
rect 8226 2313 8292 2325
<< metal2 >>
rect 4632 13533 4674 13581
rect 1791 13434 1833 13473
rect 2019 13434 2139 13473
rect 1791 13401 2139 13434
rect 2001 13368 2139 13401
rect 1923 13329 1986 13344
rect 1959 13299 1986 13329
rect 1527 13167 1686 13209
rect 1638 13143 1686 13167
rect 1638 13104 1647 13143
rect 1683 13104 1686 13143
rect 1638 12981 1686 13104
rect 1527 12861 1686 12981
rect 1923 12939 1986 13299
rect 1527 11745 1887 11790
rect 1527 10323 1842 10365
rect 1527 8901 1797 8943
rect 1527 7479 1749 7521
rect 1527 6090 1614 6093
rect 1656 6090 1701 6105
rect 1527 6054 1701 6090
rect 1551 6048 1701 6054
rect 1527 4635 1626 4683
rect 1569 4173 1626 4635
rect 1656 4242 1701 6048
rect 1716 4716 1749 7479
rect 1716 4704 1725 4716
rect 1737 4704 1749 4716
rect 1716 4701 1749 4704
rect 1764 4686 1797 8901
rect 1764 4674 1773 4686
rect 1785 4674 1797 4686
rect 1764 4671 1797 4674
rect 1809 4656 1842 10323
rect 1809 4644 1818 4656
rect 1830 4644 1842 4656
rect 1809 4641 1842 4644
rect 1854 4629 1887 11745
rect 1854 4617 1863 4629
rect 1875 4617 1887 4629
rect 1854 4614 1887 4617
rect 1926 4395 1986 12939
rect 1926 4365 1929 4395
rect 1983 4365 1986 4395
rect 1656 4212 1659 4242
rect 1695 4233 1701 4242
rect 1656 4209 1695 4212
rect 1569 4170 1641 4173
rect 1569 4131 1596 4170
rect 1569 4128 1641 4131
rect 1590 4107 1641 4113
rect 1590 4074 1602 4107
rect 1590 4068 1641 4074
rect 1590 3255 1647 4068
rect 1527 3210 1647 3255
rect 2001 2043 2061 13368
rect 3213 13329 3255 13473
rect 3213 13302 3216 13329
rect 3240 13302 3255 13329
rect 3213 13296 3255 13302
rect 2073 13251 2139 13257
rect 2073 13212 2076 13251
rect 2136 13212 2139 13251
rect 4635 13245 4677 13464
rect 7479 13389 7521 13473
rect 8901 13410 8943 13473
rect 10323 13431 10365 13473
rect 11745 13452 11787 13473
rect 11745 13440 13128 13452
rect 10323 13419 13098 13431
rect 8901 13398 13068 13410
rect 7479 13377 13035 13389
rect 4635 13218 4638 13245
rect 4662 13218 4677 13245
rect 4635 13212 4677 13218
rect 2073 13185 2139 13212
rect 2076 4791 2136 13185
rect 2076 4746 2082 4791
rect 2127 4746 2136 4791
rect 2076 4740 2136 4746
rect 2148 13143 2208 13146
rect 2148 13107 2151 13143
rect 2205 13107 2208 13143
rect 2148 2328 2208 13107
rect 10269 4839 10314 4842
rect 10269 4791 10272 4839
rect 10311 4791 10314 4839
rect 9825 4755 10104 4767
rect 9720 4737 10086 4746
rect 9720 4716 9732 4737
rect 9753 4716 10068 4728
rect 9753 4686 9765 4716
rect 9783 4698 10047 4707
rect 9783 4656 9795 4698
rect 9855 4656 9867 4659
rect 2274 4425 2286 4428
rect 4059 4353 4668 4365
rect 3447 4332 4341 4341
rect 3447 4326 3459 4332
rect 4356 4332 4383 4341
rect 3393 4314 3459 4326
rect 3393 4296 3408 4314
rect 3441 4299 3459 4314
rect 4338 4302 4359 4317
rect 3333 4287 3408 4296
rect 3441 4287 3864 4299
rect 4338 4296 4347 4302
rect 3333 4260 3357 4287
rect 3417 4272 3429 4287
rect 3468 4272 3792 4278
rect 3417 4266 3792 4272
rect 3417 4263 3618 4266
rect 3468 4260 3618 4263
rect 3492 4242 3618 4260
rect 3780 4263 3792 4266
rect 3852 4263 3864 4287
rect 4656 4284 4668 4353
rect 9855 4341 9867 4644
rect 9882 4641 9894 4644
rect 9882 4341 9894 4629
rect 9909 4626 9921 4629
rect 9909 4341 9921 4614
rect 9936 4611 9948 4614
rect 9936 4341 9948 4599
rect 5052 4305 5073 4320
rect 3300 4221 3573 4233
rect 4350 4230 4362 4251
rect 4428 4245 4437 4260
rect 5058 4242 5073 4305
rect 5103 4266 5118 4308
rect 9285 4287 9543 4296
rect 7158 4257 7200 4275
rect 9285 4257 9300 4287
rect 7158 4230 7200 4248
rect 9318 4266 9447 4278
rect 9318 4242 9333 4266
rect 9435 4248 9447 4266
rect 9531 4248 9543 4287
rect 3300 4218 3582 4221
rect 3300 4209 3576 4218
rect 7158 4203 7200 4221
rect 10038 4212 10047 4698
rect 10059 4278 10068 4716
rect 10077 4296 10086 4737
rect 10095 4356 10104 4755
rect 10269 4359 10314 4791
rect 13017 4701 13035 13377
rect 13005 4698 13035 4701
rect 13023 4689 13035 4698
rect 13050 4674 13068 13398
rect 13038 4671 13068 4674
rect 13056 4665 13068 4671
rect 13080 4647 13098 13419
rect 13071 4644 13098 4647
rect 13089 4638 13098 4644
rect 13110 4620 13128 13440
rect 13167 13344 13209 13473
rect 13104 4617 13128 4620
rect 13140 13302 13209 13344
rect 13140 4590 13155 13302
rect 13140 4566 13155 4569
rect 13173 13209 13410 13212
rect 13173 13167 13470 13209
rect 13173 13164 13410 13167
rect 13173 4545 13194 13164
rect 13203 11742 13473 11790
rect 13173 4530 13176 4545
rect 13191 4530 13194 4545
rect 13173 4527 13194 4530
rect 13206 4518 13221 11742
rect 13206 4500 13221 4503
rect 13233 10320 13473 10368
rect 13233 4491 13248 10320
rect 13260 8898 13500 8946
rect 13233 4476 13236 4491
rect 13233 4473 13248 4476
rect 13260 4461 13275 8898
rect 13272 4446 13275 4461
rect 13260 4443 13275 4446
rect 10281 4305 10335 4317
rect 10095 4263 10107 4305
rect 10323 4281 10335 4305
rect 10095 4248 10104 4263
rect 3282 4167 3366 4173
rect 3324 4161 3366 4167
rect 3357 4134 3366 4161
rect 3324 4131 3366 4134
rect 3282 4128 3366 4131
rect 3462 4104 3504 4113
rect 3495 4077 3504 4104
rect 3462 4068 3504 4077
rect 6858 3081 6951 3090
rect 6840 3051 6858 3081
rect 6951 3051 6978 3081
rect 2001 1986 2004 2043
rect 2058 1986 2061 2043
rect 2001 1983 2061 1986
rect 6018 2274 6147 2292
rect 6018 2244 6066 2274
rect 6111 2244 6147 2274
rect 3210 1965 3258 1968
rect 3210 1944 3213 1965
rect 3255 1944 3258 1965
rect 3210 1524 3258 1944
rect 4635 1923 4677 1926
rect 4635 1902 4638 1923
rect 4674 1902 4677 1923
rect 4635 1527 4677 1902
rect 6018 1566 6147 2244
rect 6840 2289 6978 3051
rect 6840 2244 6858 2289
rect 6915 2244 6978 2289
rect 6840 2229 6978 2244
rect 7008 1959 7044 3063
rect 12522 2325 12621 3063
rect 7008 1947 7011 1959
rect 7041 1947 7044 1959
rect 7458 2316 7545 2325
rect 7458 2247 7470 2316
rect 7533 2247 7545 2316
rect 6036 1563 6123 1566
rect 6054 1527 6102 1563
rect 7458 1560 7545 2247
rect 8226 2043 8292 2313
rect 12522 2241 12525 2325
rect 12618 2241 12621 2325
rect 12522 2238 12621 2241
rect 12708 2502 12744 3063
rect 8226 1986 8232 2043
rect 8286 1986 8292 2043
rect 8226 1977 8292 1986
rect 8895 2169 8934 2172
rect 8895 2151 8901 2169
rect 8895 1914 8934 2151
rect 10323 2127 10362 2130
rect 10323 2106 10329 2127
rect 10359 2106 10362 2127
rect 7479 1527 7521 1560
rect 8892 1551 8940 1914
rect 10323 1899 10362 2106
rect 11754 1923 11784 2064
rect 12708 1923 12747 2502
rect 13194 2196 13197 2217
rect 13176 1947 13197 2196
rect 8895 1527 8940 1551
rect 10317 1527 10365 1899
rect 11742 1527 11790 1923
rect 12708 1902 12711 1923
rect 12744 1902 12747 1923
rect 12708 1899 12747 1902
rect 13164 1527 13212 1947
<< m3contact >>
rect 1923 13299 1959 13329
rect 1647 13104 1683 13143
rect 1725 4704 1737 4716
rect 1773 4674 1785 4686
rect 1818 4644 1830 4656
rect 1863 4617 1875 4629
rect 1929 4356 1983 4395
rect 1659 4212 1695 4242
rect 1596 4131 1641 4170
rect 1602 4074 1641 4107
rect 3216 13302 3240 13329
rect 2076 13212 2136 13251
rect 4638 13218 4662 13245
rect 2082 4746 2127 4791
rect 2151 13107 2205 13143
rect 10272 4791 10311 4839
rect 9813 4755 9825 4767
rect 9720 4704 9732 4716
rect 9753 4674 9765 4686
rect 9783 4644 9795 4656
rect 9855 4644 9867 4656
rect 9813 4617 9825 4629
rect 7893 4587 7908 4602
rect 2274 4428 2289 4443
rect 4032 4353 4059 4380
rect 4341 4329 4356 4344
rect 4410 4320 4425 4335
rect 4590 4305 4605 4320
rect 4347 4287 4362 4302
rect 4380 4269 4395 4287
rect 9855 4329 9867 4341
rect 9882 4629 9894 4641
rect 9882 4329 9894 4341
rect 9909 4614 9921 4626
rect 9909 4329 9921 4341
rect 9936 4599 9948 4611
rect 9936 4329 9948 4341
rect 5037 4305 5052 4320
rect 3270 4209 3300 4233
rect 4437 4245 4452 4260
rect 5103 4308 5118 4323
rect 13005 4680 13023 4698
rect 13038 4653 13056 4671
rect 13071 4626 13089 4644
rect 13104 4599 13122 4617
rect 13137 4569 13155 4590
rect 13176 4530 13191 4545
rect 13206 4503 13221 4518
rect 13236 4476 13251 4491
rect 13257 4446 13272 4461
rect 3282 4131 3324 4167
rect 4188 4116 4203 4131
rect 9855 4113 9870 4128
rect 4188 4044 4203 4059
rect 9855 4041 9870 4056
rect 4188 3972 4203 3987
rect 9855 3969 9870 3984
rect 4188 3900 4203 3915
rect 9855 3897 9870 3912
rect 2004 1986 2058 2043
rect 6066 2244 6111 2274
rect 3213 1944 3255 1965
rect 4638 1902 4674 1923
rect 6858 2244 6915 2289
rect 7011 1947 7041 1959
rect 7470 2247 7533 2316
rect 12525 2241 12618 2325
rect 8232 1986 8286 2043
rect 8901 2151 8934 2169
rect 10329 2106 10359 2127
rect 11748 2064 11784 2082
rect 13173 2196 13194 2217
rect 12711 1902 12744 1923
<< metal3 >>
rect 1914 13329 3261 13341
rect 1914 13299 1923 13329
rect 1959 13302 3216 13329
rect 3240 13302 3261 13329
rect 1959 13299 3261 13302
rect 1914 13290 3261 13299
rect 2073 13251 4683 13257
rect 2073 13212 2076 13251
rect 2136 13245 4683 13251
rect 2136 13218 4638 13245
rect 4662 13218 4683 13245
rect 2136 13212 4683 13218
rect 2073 13206 4683 13212
rect 1641 13143 2208 13149
rect 1641 13104 1647 13143
rect 1683 13107 2151 13143
rect 2205 13107 2208 13143
rect 1683 13104 2208 13107
rect 1641 13098 2208 13104
rect 9612 4839 10314 4842
rect 9612 4797 10272 4839
rect 2076 4791 10272 4797
rect 10311 4791 10314 4839
rect 2076 4746 2082 4791
rect 2127 4788 10314 4791
rect 2127 4746 9654 4788
rect 2076 4740 9654 4746
rect 9810 4767 9828 4770
rect 9810 4755 9813 4767
rect 9825 4755 9828 4767
rect 1722 4716 9735 4719
rect 1722 4704 1725 4716
rect 1737 4704 9720 4716
rect 9732 4704 9735 4716
rect 1722 4701 9735 4704
rect 1770 4686 9768 4689
rect 1770 4674 1773 4686
rect 1785 4674 9753 4686
rect 9765 4674 9768 4686
rect 1770 4671 9768 4674
rect 1815 4656 9798 4659
rect 1815 4644 1818 4656
rect 1830 4644 9783 4656
rect 9795 4644 9798 4656
rect 1815 4641 9798 4644
rect 9810 4632 9828 4755
rect 13002 4698 13026 4701
rect 13002 4686 13005 4698
rect 9852 4680 13005 4686
rect 13023 4680 13026 4698
rect 9852 4671 13026 4680
rect 13035 4671 13059 4674
rect 9852 4656 9870 4671
rect 13035 4662 13038 4671
rect 9852 4644 9855 4656
rect 9867 4644 9870 4656
rect 9852 4641 9870 4644
rect 9879 4653 13038 4662
rect 13056 4653 13059 4671
rect 9879 4647 13059 4653
rect 9879 4641 9897 4647
rect 1860 4629 9828 4632
rect 1860 4617 1863 4629
rect 1875 4617 9813 4629
rect 9825 4617 9828 4629
rect 9879 4629 9882 4641
rect 9894 4629 9897 4641
rect 13068 4644 13092 4647
rect 13068 4638 13071 4644
rect 9879 4626 9897 4629
rect 9906 4626 13071 4638
rect 13089 4626 13092 4644
rect 1860 4614 9828 4617
rect 9906 4614 9909 4626
rect 9921 4623 13092 4626
rect 9921 4614 9924 4623
rect 13101 4617 13125 4620
rect 9906 4611 9924 4614
rect 9933 4611 9951 4614
rect 13101 4611 13104 4617
rect 7890 4602 7911 4605
rect 7890 4587 7893 4602
rect 7908 4587 7911 4602
rect 9933 4599 9936 4611
rect 9948 4599 13104 4611
rect 13122 4599 13125 4617
rect 9933 4596 13125 4599
rect 13134 4590 13158 4593
rect 13134 4587 13137 4590
rect 2214 4569 13137 4587
rect 13155 4569 13158 4590
rect 2217 4467 2232 4569
rect 13134 4566 13158 4569
rect 13173 4545 13194 4548
rect 4191 4530 13176 4545
rect 13191 4530 13194 4545
rect 4191 4527 13194 4530
rect 2217 4452 2292 4467
rect 2271 4443 2292 4452
rect 2271 4428 2274 4443
rect 2289 4428 2292 4443
rect 2271 4425 2292 4428
rect 1926 4395 2010 4398
rect 1926 4356 1929 4395
rect 1983 4383 2010 4395
rect 1983 4380 4062 4383
rect 1983 4356 4032 4380
rect 1926 4353 4032 4356
rect 4059 4353 4062 4380
rect 4029 4350 4062 4353
rect 1656 4242 1701 4245
rect 1656 4212 1659 4242
rect 1695 4236 1701 4242
rect 1695 4233 3303 4236
rect 1695 4212 3270 4233
rect 1656 4209 3270 4212
rect 3300 4209 3303 4233
rect 3267 4206 3303 4209
rect 1593 4170 3333 4173
rect 1593 4131 1596 4170
rect 1641 4167 3333 4170
rect 1641 4131 3282 4167
rect 3324 4131 3333 4167
rect 4191 4134 4206 4527
rect 13203 4518 13224 4521
rect 1593 4128 3333 4131
rect 4185 4131 4206 4134
rect 4185 4116 4188 4131
rect 4203 4116 4206 4131
rect 4185 4113 4206 4116
rect 4215 4503 13206 4518
rect 13221 4503 13224 4518
rect 4215 4500 13224 4503
rect 1590 4107 3465 4113
rect 1590 4074 1602 4107
rect 1641 4074 3465 4107
rect 1590 4068 3465 4074
rect 4185 4059 4206 4062
rect 4185 4044 4188 4059
rect 4203 4056 4206 4059
rect 4215 4056 4230 4500
rect 13233 4491 13254 4494
rect 4203 4044 4230 4056
rect 4185 4041 4230 4044
rect 4239 4476 13236 4491
rect 13251 4476 13254 4491
rect 4239 4473 13254 4476
rect 4185 3987 4206 3990
rect 4185 3972 4188 3987
rect 4203 3984 4206 3987
rect 4239 3984 4254 4473
rect 4203 3972 4254 3984
rect 4185 3969 4254 3972
rect 4263 4461 13275 4464
rect 4263 4446 13257 4461
rect 13272 4446 13275 4461
rect 4185 3915 4206 3918
rect 4185 3900 4188 3915
rect 4203 3912 4206 3915
rect 4263 3912 4278 4446
rect 13254 4443 13275 4446
rect 4338 4347 5121 4362
rect 4338 4344 4359 4347
rect 4338 4329 4341 4344
rect 4356 4329 4359 4344
rect 4338 4326 4359 4329
rect 4407 4335 4428 4338
rect 4407 4320 4410 4335
rect 4425 4320 4428 4335
rect 5100 4323 5121 4347
rect 9852 4341 9870 4344
rect 9852 4329 9855 4341
rect 9867 4329 9870 4341
rect 9852 4326 9870 4329
rect 9879 4341 9897 4344
rect 9879 4329 9882 4341
rect 9894 4329 9897 4341
rect 9879 4326 9897 4329
rect 4407 4317 4428 4320
rect 4587 4320 5055 4323
rect 4344 4302 4365 4305
rect 4344 4287 4347 4302
rect 4362 4287 4365 4302
rect 4344 4239 4365 4287
rect 4377 4287 4398 4290
rect 4377 4269 4380 4287
rect 4395 4269 4398 4287
rect 4377 4266 4398 4269
rect 4203 3900 4302 3912
rect 4185 3897 4302 3900
rect 4350 2133 4365 4239
rect 4347 2088 4365 2133
rect 4383 2130 4398 4266
rect 4407 2172 4422 4317
rect 4587 4305 4590 4320
rect 4605 4305 5037 4320
rect 5052 4305 5055 4320
rect 5100 4308 5103 4323
rect 5118 4308 5121 4323
rect 5100 4305 5121 4308
rect 9855 4317 9870 4326
rect 4587 4302 5055 4305
rect 9855 4299 9873 4317
rect 4434 4260 4455 4263
rect 4431 4245 4437 4260
rect 4452 4245 4455 4260
rect 4431 4242 4455 4245
rect 4431 4239 4452 4242
rect 4431 2220 4446 4239
rect 9858 4131 9873 4299
rect 9852 4128 9873 4131
rect 9852 4113 9855 4128
rect 9870 4113 9873 4128
rect 9852 4110 9873 4113
rect 9882 4059 9897 4326
rect 9852 4056 9897 4059
rect 9852 4041 9855 4056
rect 9870 4041 9897 4056
rect 9852 4038 9897 4041
rect 9906 4341 9924 4344
rect 9906 4329 9909 4341
rect 9921 4329 9924 4341
rect 9906 4326 9924 4329
rect 9933 4341 9951 4344
rect 9933 4329 9936 4341
rect 9948 4329 9951 4341
rect 9933 4326 9951 4329
rect 9906 3987 9921 4326
rect 9933 4317 9948 4326
rect 9852 3984 9921 3987
rect 9852 3969 9855 3984
rect 9870 3969 9921 3984
rect 9852 3966 9921 3969
rect 9930 4302 9948 4317
rect 9930 3915 9945 4302
rect 9852 3912 9945 3915
rect 9852 3897 9855 3912
rect 9870 3897 9945 3912
rect 9852 3894 9945 3897
rect 6051 2289 6933 2361
rect 6051 2274 6858 2289
rect 6051 2244 6066 2274
rect 6111 2244 6858 2274
rect 6915 2244 6933 2289
rect 6051 2229 6933 2244
rect 7458 2325 12621 2328
rect 7458 2316 12525 2325
rect 7458 2247 7470 2316
rect 7533 2247 12525 2316
rect 7458 2241 12525 2247
rect 12618 2241 12621 2325
rect 7458 2238 12621 2241
rect 4431 2217 13197 2220
rect 4431 2196 13173 2217
rect 13194 2196 13197 2217
rect 4431 2193 13197 2196
rect 4407 2169 8937 2172
rect 4407 2151 8901 2169
rect 8934 2151 8937 2169
rect 4407 2145 8937 2151
rect 4383 2127 10362 2130
rect 4383 2106 10329 2127
rect 10359 2106 10362 2127
rect 4383 2103 10362 2106
rect 4347 2082 11787 2088
rect 4347 2064 11748 2082
rect 11784 2064 11787 2082
rect 4347 2061 11787 2064
rect 2001 2043 8289 2046
rect 2001 1986 2004 2043
rect 2058 1986 8232 2043
rect 8286 1986 8289 2043
rect 2001 1983 8289 1986
rect 3210 1965 7044 1968
rect 3210 1944 3213 1965
rect 3255 1959 7044 1965
rect 3255 1947 7011 1959
rect 7041 1947 7044 1959
rect 3255 1944 7044 1947
rect 3210 1941 7044 1944
rect 4635 1923 12747 1926
rect 4635 1902 4638 1923
rect 4674 1902 12711 1923
rect 12744 1902 12747 1923
rect 4635 1899 12747 1902
use barepad  barepad_1
timestamp 1259953556
transform -1 0 2523 0 -1 15000
box -6 0 1428 1539
use inpad  inpad_1
timestamp 1259953556
transform -1 0 3945 0 -1 15000
box -6 0 1428 1539
use inpad  inpad_0
timestamp 1259953556
transform -1 0 5367 0 -1 15000
box -6 0 1428 1539
use blankpad  blankpad_3
timestamp 1259953556
transform -1 0 6789 0 -1 15000
box -6 0 1428 1539
use inorpad  inorpad_6
timestamp 1259953556
transform -1 0 8211 0 -1 15000
box -6 0 1428 1539
use inorpad  inorpad_5
timestamp 1259953556
transform -1 0 9633 0 -1 15000
box -6 0 1428 1539
use inorpad  inorpad_4
timestamp 1259953556
transform -1 0 11055 0 -1 15000
box -6 0 1428 1539
use inorpad  inorpad_3
timestamp 1259953556
transform -1 0 12477 0 -1 15000
box -6 0 1428 1539
use barepad  barepad_0
timestamp 1259953556
transform -1 0 13899 0 -1 15000
box -6 0 1428 1539
use padframe_top  padframe_top_0
timestamp 1259953556
transform 1 0 0 0 1 13461
box 0 0 15000 1539
use barepad  barepad_2
timestamp 1259953556
transform 0 1 0 -1 0 13899
box -6 0 1428 1539
use inorpad  inorpad_17
timestamp 1259953556
transform 0 -1 15000 1 0 12477
box -6 0 1428 1539
use inorpad  inorpad_7
timestamp 1259953556
transform 0 1 0 -1 0 12477
box -6 0 1428 1539
use inorpad  inorpad_8
timestamp 1259953556
transform 0 1 0 -1 0 11055
box -6 0 1428 1539
use inorpad  inorpad_9
timestamp 1259953556
transform 0 1 0 -1 0 9633
box -6 0 1428 1539
use inorpad  inorpad_10
timestamp 1259953556
transform 0 1 0 -1 0 8211
box -6 0 1428 1539
use inpad  inpad_2
timestamp 1259953556
transform 0 1 0 -1 0 6789
box -6 0 1428 1539
use forrest-threshold  forrest-threshold_0
timestamp 1419146600
transform 1 0 2226 0 1 4770
box 45 78 10691 7457
use inorpad  inorpad_0
timestamp 1259953556
transform 0 -1 15000 1 0 11055
box -6 0 1428 1539
use inorpad  inorpad_1
timestamp 1259953556
transform 0 -1 15000 1 0 9633
box -6 0 1428 1539
use inorpad  inorpad_2
timestamp 1259953556
transform 0 -1 15000 1 0 8211
box -6 0 1428 1539
use blankpad  blankpad_2
timestamp 1259953556
transform 0 -1 15000 1 0 6789
box -6 0 1428 1539
use blankpad  blankpad_7
timestamp 1259953556
transform 0 -1 15000 1 0 5367
box -6 0 1428 1539
use inpad  inpad_3
timestamp 1259953556
transform 0 1 0 -1 0 5367
box -6 0 1428 1539
use inpad  inpad_4
timestamp 1259953556
transform 0 1 0 -1 0 3945
box -6 0 1428 1539
use top-level  top-level_0
timestamp 1419034691
transform 1 0 2115 0 1 2316
box 0 0 5199 2133
use top-level  top-level_1
timestamp 1419034691
transform 1 0 7782 0 1 2313
box 0 0 5199 2133
use blankpad  blankpad_8
timestamp 1259953556
transform 0 -1 15000 1 0 3945
box -6 0 1428 1539
use blankpad  blankpad_1
timestamp 1259953556
transform 0 -1 15000 1 0 2523
box -6 0 1428 1539
use padframe_left  padframe_left_0
timestamp 1259953556
transform 1 0 0 0 1 1101
box 6 6 1539 12792
use barepad  barepad_4
timestamp 1259953556
transform 0 1 0 -1 0 2523
box -6 0 1428 1539
use barepad  barepad_3
timestamp 1259953556
transform 1 0 1101 0 1 0
box -6 0 1428 1539
use inorpad  inorpad_11
timestamp 1259953556
transform 1 0 2523 0 1 0
box -6 0 1428 1539
use inorpad  inorpad_12
timestamp 1259953556
transform 1 0 3945 0 1 0
box -6 0 1428 1539
use inorpad  inorpad_18
timestamp 1259953556
transform 1 0 5367 0 1 0
box -6 0 1428 1539
use inorpad  inorpad_19
timestamp 1259953556
transform 1 0 6789 0 1 0
box -6 0 1428 1539
use inorpad  inorpad_13
timestamp 1259953556
transform 1 0 8211 0 1 0
box -6 0 1428 1539
use inorpad  inorpad_14
timestamp 1259953556
transform 1 0 9633 0 1 0
box -6 0 1428 1539
use inorpad  inorpad_15
timestamp 1259953556
transform 1 0 11055 0 1 0
box -6 0 1428 1539
use padframe_right  padframe_right_0
timestamp 1259953556
transform 1 0 13461 0 1 1101
box 0 6 1533 12792
use blankpad  blankpad_0
timestamp 1259953556
transform 0 -1 15000 1 0 1101
box -6 0 1428 1539
use inorpad  inorpad_16
timestamp 1259953556
transform 1 0 12477 0 1 0
box -6 0 1428 1539
use padframe_bottom  padframe_bottom_0
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 15000 1539
<< labels >>
rlabel space 4188 4245 4206 4254 1 x1
rlabel space 4212 4245 4230 4254 1 x2
rlabel space 4236 4245 4254 4254 1 x3
rlabel space 4260 4245 4278 4254 1 x4
rlabel metal3 9858 4248 9873 4254 1 x1
rlabel metal3 9882 4248 9897 4254 1 x2
rlabel metal3 9906 4248 9921 4254 1 x3
rlabel metal3 9930 4248 9945 4254 1 x4
rlabel metal3 9777 4614 9825 4632 1 20
rlabel metal3 9717 4671 9765 4689 1 18
rlabel metal3 9747 4641 9795 4659 1 19
rlabel metal3 9687 4701 9735 4719 1 17
<< end >>
