magic
tech scmos
timestamp 1259953556
<< electrodecontact >>
rect 539 489 543 493
rect 545 489 549 493
rect 551 489 555 493
rect 557 489 561 493
rect 563 489 567 493
rect 569 489 573 493
rect 575 489 579 493
rect 539 471 543 475
rect 545 471 549 475
rect 551 471 555 475
rect 557 471 561 475
rect 563 471 567 475
rect 569 471 573 475
rect 575 471 579 475
rect 573 456 577 460
rect 583 456 587 460
rect 629 489 633 493
rect 635 489 639 493
rect 641 489 645 493
rect 647 489 651 493
rect 653 489 657 493
rect 659 489 663 493
rect 665 489 669 493
rect 629 471 633 475
rect 635 471 639 475
rect 641 471 645 475
rect 647 471 651 475
rect 653 471 657 475
rect 659 471 663 475
rect 665 471 669 475
rect 621 456 625 460
rect 631 456 635 460
rect 540 445 544 449
rect 546 445 550 449
rect 552 445 556 449
rect 558 445 562 449
rect 564 445 568 449
rect 540 439 544 443
rect 546 439 550 443
rect 552 439 556 443
rect 558 439 562 443
rect 564 439 568 443
rect 540 433 544 437
rect 546 433 550 437
rect 552 433 556 437
rect 558 433 562 437
rect 564 433 568 437
rect 540 427 544 431
rect 546 427 550 431
rect 552 427 556 431
rect 558 427 562 431
rect 564 427 568 431
rect 540 420 544 424
rect 546 420 550 424
rect 552 420 556 424
rect 558 420 562 424
rect 564 420 568 424
rect 540 414 544 418
rect 546 414 550 418
rect 552 414 556 418
rect 558 414 562 418
rect 564 414 568 418
rect 640 445 644 449
rect 646 445 650 449
rect 652 445 656 449
rect 658 445 662 449
rect 664 445 668 449
rect 640 439 644 443
rect 646 439 650 443
rect 652 439 656 443
rect 658 439 662 443
rect 664 439 668 443
rect 640 433 644 437
rect 646 433 650 437
rect 652 433 656 437
rect 658 433 662 437
rect 664 433 668 437
rect 640 427 644 431
rect 646 427 650 431
rect 652 427 656 431
rect 658 427 662 431
rect 664 427 668 431
rect 640 420 644 424
rect 646 420 650 424
rect 652 420 656 424
rect 658 420 662 424
rect 664 420 668 424
rect 640 414 644 418
rect 646 414 650 418
rect 652 414 656 418
rect 658 414 662 418
rect 664 414 668 418
rect 539 397 543 401
rect 545 397 549 401
rect 551 397 555 401
rect 557 397 561 401
rect 563 397 567 401
rect 569 397 573 401
rect 575 397 579 401
rect 539 384 543 388
rect 545 384 549 388
rect 551 384 555 388
rect 557 384 561 388
rect 563 384 567 388
rect 569 384 573 388
rect 575 384 579 388
rect 629 397 633 401
rect 635 397 639 401
rect 641 397 645 401
rect 647 397 651 401
rect 653 397 657 401
rect 659 397 663 401
rect 665 397 669 401
rect 629 384 633 388
rect 635 384 639 388
rect 641 384 645 388
rect 647 384 651 388
rect 653 384 657 388
rect 659 384 663 388
rect 665 384 669 388
rect 1013 489 1017 493
rect 1019 489 1023 493
rect 1025 489 1029 493
rect 1031 489 1035 493
rect 1037 489 1041 493
rect 1043 489 1047 493
rect 1049 489 1053 493
rect 1013 471 1017 475
rect 1019 471 1023 475
rect 1025 471 1029 475
rect 1031 471 1035 475
rect 1037 471 1041 475
rect 1043 471 1047 475
rect 1049 471 1053 475
rect 1047 456 1051 460
rect 1057 456 1061 460
rect 1103 489 1107 493
rect 1109 489 1113 493
rect 1115 489 1119 493
rect 1121 489 1125 493
rect 1127 489 1131 493
rect 1133 489 1137 493
rect 1139 489 1143 493
rect 1103 471 1107 475
rect 1109 471 1113 475
rect 1115 471 1119 475
rect 1121 471 1125 475
rect 1127 471 1131 475
rect 1133 471 1137 475
rect 1139 471 1143 475
rect 1095 456 1099 460
rect 1105 456 1109 460
rect 1014 445 1018 449
rect 1020 445 1024 449
rect 1026 445 1030 449
rect 1032 445 1036 449
rect 1038 445 1042 449
rect 1014 439 1018 443
rect 1020 439 1024 443
rect 1026 439 1030 443
rect 1032 439 1036 443
rect 1038 439 1042 443
rect 1014 433 1018 437
rect 1020 433 1024 437
rect 1026 433 1030 437
rect 1032 433 1036 437
rect 1038 433 1042 437
rect 1014 427 1018 431
rect 1020 427 1024 431
rect 1026 427 1030 431
rect 1032 427 1036 431
rect 1038 427 1042 431
rect 1014 420 1018 424
rect 1020 420 1024 424
rect 1026 420 1030 424
rect 1032 420 1036 424
rect 1038 420 1042 424
rect 1014 414 1018 418
rect 1020 414 1024 418
rect 1026 414 1030 418
rect 1032 414 1036 418
rect 1038 414 1042 418
rect 1114 445 1118 449
rect 1120 445 1124 449
rect 1126 445 1130 449
rect 1132 445 1136 449
rect 1138 445 1142 449
rect 1114 439 1118 443
rect 1120 439 1124 443
rect 1126 439 1130 443
rect 1132 439 1136 443
rect 1138 439 1142 443
rect 1114 433 1118 437
rect 1120 433 1124 437
rect 1126 433 1130 437
rect 1132 433 1136 437
rect 1138 433 1142 437
rect 1114 427 1118 431
rect 1120 427 1124 431
rect 1126 427 1130 431
rect 1132 427 1136 431
rect 1138 427 1142 431
rect 1114 420 1118 424
rect 1120 420 1124 424
rect 1126 420 1130 424
rect 1132 420 1136 424
rect 1138 420 1142 424
rect 1114 414 1118 418
rect 1120 414 1124 418
rect 1126 414 1130 418
rect 1132 414 1136 418
rect 1138 414 1142 418
rect 1013 397 1017 401
rect 1019 397 1023 401
rect 1025 397 1029 401
rect 1031 397 1035 401
rect 1037 397 1041 401
rect 1043 397 1047 401
rect 1049 397 1053 401
rect 1013 384 1017 388
rect 1019 384 1023 388
rect 1025 384 1029 388
rect 1031 384 1035 388
rect 1037 384 1041 388
rect 1043 384 1047 388
rect 1049 384 1053 388
rect 1103 397 1107 401
rect 1109 397 1113 401
rect 1115 397 1119 401
rect 1121 397 1125 401
rect 1127 397 1131 401
rect 1133 397 1137 401
rect 1139 397 1143 401
rect 1103 384 1107 388
rect 1109 384 1113 388
rect 1115 384 1119 388
rect 1121 384 1125 388
rect 1127 384 1131 388
rect 1133 384 1137 388
rect 1139 384 1143 388
rect 1487 489 1491 493
rect 1493 489 1497 493
rect 1499 489 1503 493
rect 1505 489 1509 493
rect 1511 489 1515 493
rect 1517 489 1521 493
rect 1523 489 1527 493
rect 1487 471 1491 475
rect 1493 471 1497 475
rect 1499 471 1503 475
rect 1505 471 1509 475
rect 1511 471 1515 475
rect 1517 471 1521 475
rect 1523 471 1527 475
rect 1521 456 1525 460
rect 1531 456 1535 460
rect 1577 489 1581 493
rect 1583 489 1587 493
rect 1589 489 1593 493
rect 1595 489 1599 493
rect 1601 489 1605 493
rect 1607 489 1611 493
rect 1613 489 1617 493
rect 1577 471 1581 475
rect 1583 471 1587 475
rect 1589 471 1593 475
rect 1595 471 1599 475
rect 1601 471 1605 475
rect 1607 471 1611 475
rect 1613 471 1617 475
rect 1569 456 1573 460
rect 1579 456 1583 460
rect 1488 445 1492 449
rect 1494 445 1498 449
rect 1500 445 1504 449
rect 1506 445 1510 449
rect 1512 445 1516 449
rect 1488 439 1492 443
rect 1494 439 1498 443
rect 1500 439 1504 443
rect 1506 439 1510 443
rect 1512 439 1516 443
rect 1488 433 1492 437
rect 1494 433 1498 437
rect 1500 433 1504 437
rect 1506 433 1510 437
rect 1512 433 1516 437
rect 1488 427 1492 431
rect 1494 427 1498 431
rect 1500 427 1504 431
rect 1506 427 1510 431
rect 1512 427 1516 431
rect 1488 420 1492 424
rect 1494 420 1498 424
rect 1500 420 1504 424
rect 1506 420 1510 424
rect 1512 420 1516 424
rect 1488 414 1492 418
rect 1494 414 1498 418
rect 1500 414 1504 418
rect 1506 414 1510 418
rect 1512 414 1516 418
rect 1588 445 1592 449
rect 1594 445 1598 449
rect 1600 445 1604 449
rect 1606 445 1610 449
rect 1612 445 1616 449
rect 1588 439 1592 443
rect 1594 439 1598 443
rect 1600 439 1604 443
rect 1606 439 1610 443
rect 1612 439 1616 443
rect 1588 433 1592 437
rect 1594 433 1598 437
rect 1600 433 1604 437
rect 1606 433 1610 437
rect 1612 433 1616 437
rect 1588 427 1592 431
rect 1594 427 1598 431
rect 1600 427 1604 431
rect 1606 427 1610 431
rect 1612 427 1616 431
rect 1588 420 1592 424
rect 1594 420 1598 424
rect 1600 420 1604 424
rect 1606 420 1610 424
rect 1612 420 1616 424
rect 1588 414 1592 418
rect 1594 414 1598 418
rect 1600 414 1604 418
rect 1606 414 1610 418
rect 1612 414 1616 418
rect 1487 397 1491 401
rect 1493 397 1497 401
rect 1499 397 1503 401
rect 1505 397 1509 401
rect 1511 397 1515 401
rect 1517 397 1521 401
rect 1523 397 1527 401
rect 1487 384 1491 388
rect 1493 384 1497 388
rect 1499 384 1503 388
rect 1505 384 1509 388
rect 1511 384 1515 388
rect 1517 384 1521 388
rect 1523 384 1527 388
rect 1577 397 1581 401
rect 1583 397 1587 401
rect 1589 397 1593 401
rect 1595 397 1599 401
rect 1601 397 1605 401
rect 1607 397 1611 401
rect 1613 397 1617 401
rect 1577 384 1581 388
rect 1583 384 1587 388
rect 1589 384 1593 388
rect 1595 384 1599 388
rect 1601 384 1605 388
rect 1607 384 1611 388
rect 1613 384 1617 388
rect 1961 489 1965 493
rect 1967 489 1971 493
rect 1973 489 1977 493
rect 1979 489 1983 493
rect 1985 489 1989 493
rect 1991 489 1995 493
rect 1997 489 2001 493
rect 1961 471 1965 475
rect 1967 471 1971 475
rect 1973 471 1977 475
rect 1979 471 1983 475
rect 1985 471 1989 475
rect 1991 471 1995 475
rect 1997 471 2001 475
rect 1995 456 1999 460
rect 2005 456 2009 460
rect 2051 489 2055 493
rect 2057 489 2061 493
rect 2063 489 2067 493
rect 2069 489 2073 493
rect 2075 489 2079 493
rect 2081 489 2085 493
rect 2087 489 2091 493
rect 2051 471 2055 475
rect 2057 471 2061 475
rect 2063 471 2067 475
rect 2069 471 2073 475
rect 2075 471 2079 475
rect 2081 471 2085 475
rect 2087 471 2091 475
rect 2043 456 2047 460
rect 2053 456 2057 460
rect 1962 445 1966 449
rect 1968 445 1972 449
rect 1974 445 1978 449
rect 1980 445 1984 449
rect 1986 445 1990 449
rect 1962 439 1966 443
rect 1968 439 1972 443
rect 1974 439 1978 443
rect 1980 439 1984 443
rect 1986 439 1990 443
rect 1962 433 1966 437
rect 1968 433 1972 437
rect 1974 433 1978 437
rect 1980 433 1984 437
rect 1986 433 1990 437
rect 1962 427 1966 431
rect 1968 427 1972 431
rect 1974 427 1978 431
rect 1980 427 1984 431
rect 1986 427 1990 431
rect 1962 420 1966 424
rect 1968 420 1972 424
rect 1974 420 1978 424
rect 1980 420 1984 424
rect 1986 420 1990 424
rect 1962 414 1966 418
rect 1968 414 1972 418
rect 1974 414 1978 418
rect 1980 414 1984 418
rect 1986 414 1990 418
rect 2062 445 2066 449
rect 2068 445 2072 449
rect 2074 445 2078 449
rect 2080 445 2084 449
rect 2086 445 2090 449
rect 2062 439 2066 443
rect 2068 439 2072 443
rect 2074 439 2078 443
rect 2080 439 2084 443
rect 2086 439 2090 443
rect 2062 433 2066 437
rect 2068 433 2072 437
rect 2074 433 2078 437
rect 2080 433 2084 437
rect 2086 433 2090 437
rect 2062 427 2066 431
rect 2068 427 2072 431
rect 2074 427 2078 431
rect 2080 427 2084 431
rect 2086 427 2090 431
rect 2062 420 2066 424
rect 2068 420 2072 424
rect 2074 420 2078 424
rect 2080 420 2084 424
rect 2086 420 2090 424
rect 2062 414 2066 418
rect 2068 414 2072 418
rect 2074 414 2078 418
rect 2080 414 2084 418
rect 2086 414 2090 418
rect 1961 397 1965 401
rect 1967 397 1971 401
rect 1973 397 1977 401
rect 1979 397 1983 401
rect 1985 397 1989 401
rect 1991 397 1995 401
rect 1997 397 2001 401
rect 1961 384 1965 388
rect 1967 384 1971 388
rect 1973 384 1977 388
rect 1979 384 1983 388
rect 1985 384 1989 388
rect 1991 384 1995 388
rect 1997 384 2001 388
rect 2051 397 2055 401
rect 2057 397 2061 401
rect 2063 397 2067 401
rect 2069 397 2073 401
rect 2075 397 2079 401
rect 2081 397 2085 401
rect 2087 397 2091 401
rect 2051 384 2055 388
rect 2057 384 2061 388
rect 2063 384 2067 388
rect 2069 384 2073 388
rect 2075 384 2079 388
rect 2081 384 2085 388
rect 2087 384 2091 388
rect 2435 489 2439 493
rect 2441 489 2445 493
rect 2447 489 2451 493
rect 2453 489 2457 493
rect 2459 489 2463 493
rect 2465 489 2469 493
rect 2471 489 2475 493
rect 2435 471 2439 475
rect 2441 471 2445 475
rect 2447 471 2451 475
rect 2453 471 2457 475
rect 2459 471 2463 475
rect 2465 471 2469 475
rect 2471 471 2475 475
rect 2469 456 2473 460
rect 2479 456 2483 460
rect 2525 489 2529 493
rect 2531 489 2535 493
rect 2537 489 2541 493
rect 2543 489 2547 493
rect 2549 489 2553 493
rect 2555 489 2559 493
rect 2561 489 2565 493
rect 2525 471 2529 475
rect 2531 471 2535 475
rect 2537 471 2541 475
rect 2543 471 2547 475
rect 2549 471 2553 475
rect 2555 471 2559 475
rect 2561 471 2565 475
rect 2517 456 2521 460
rect 2527 456 2531 460
rect 2436 445 2440 449
rect 2442 445 2446 449
rect 2448 445 2452 449
rect 2454 445 2458 449
rect 2460 445 2464 449
rect 2436 439 2440 443
rect 2442 439 2446 443
rect 2448 439 2452 443
rect 2454 439 2458 443
rect 2460 439 2464 443
rect 2436 433 2440 437
rect 2442 433 2446 437
rect 2448 433 2452 437
rect 2454 433 2458 437
rect 2460 433 2464 437
rect 2436 427 2440 431
rect 2442 427 2446 431
rect 2448 427 2452 431
rect 2454 427 2458 431
rect 2460 427 2464 431
rect 2436 420 2440 424
rect 2442 420 2446 424
rect 2448 420 2452 424
rect 2454 420 2458 424
rect 2460 420 2464 424
rect 2436 414 2440 418
rect 2442 414 2446 418
rect 2448 414 2452 418
rect 2454 414 2458 418
rect 2460 414 2464 418
rect 2536 445 2540 449
rect 2542 445 2546 449
rect 2548 445 2552 449
rect 2554 445 2558 449
rect 2560 445 2564 449
rect 2536 439 2540 443
rect 2542 439 2546 443
rect 2548 439 2552 443
rect 2554 439 2558 443
rect 2560 439 2564 443
rect 2536 433 2540 437
rect 2542 433 2546 437
rect 2548 433 2552 437
rect 2554 433 2558 437
rect 2560 433 2564 437
rect 2536 427 2540 431
rect 2542 427 2546 431
rect 2548 427 2552 431
rect 2554 427 2558 431
rect 2560 427 2564 431
rect 2536 420 2540 424
rect 2542 420 2546 424
rect 2548 420 2552 424
rect 2554 420 2558 424
rect 2560 420 2564 424
rect 2536 414 2540 418
rect 2542 414 2546 418
rect 2548 414 2552 418
rect 2554 414 2558 418
rect 2560 414 2564 418
rect 2435 397 2439 401
rect 2441 397 2445 401
rect 2447 397 2451 401
rect 2453 397 2457 401
rect 2459 397 2463 401
rect 2465 397 2469 401
rect 2471 397 2475 401
rect 2435 384 2439 388
rect 2441 384 2445 388
rect 2447 384 2451 388
rect 2453 384 2457 388
rect 2459 384 2463 388
rect 2465 384 2469 388
rect 2471 384 2475 388
rect 2525 397 2529 401
rect 2531 397 2535 401
rect 2537 397 2541 401
rect 2543 397 2547 401
rect 2549 397 2553 401
rect 2555 397 2559 401
rect 2561 397 2565 401
rect 2525 384 2529 388
rect 2531 384 2535 388
rect 2537 384 2541 388
rect 2543 384 2547 388
rect 2549 384 2553 388
rect 2555 384 2559 388
rect 2561 384 2565 388
rect 2909 489 2913 493
rect 2915 489 2919 493
rect 2921 489 2925 493
rect 2927 489 2931 493
rect 2933 489 2937 493
rect 2939 489 2943 493
rect 2945 489 2949 493
rect 2909 471 2913 475
rect 2915 471 2919 475
rect 2921 471 2925 475
rect 2927 471 2931 475
rect 2933 471 2937 475
rect 2939 471 2943 475
rect 2945 471 2949 475
rect 2943 456 2947 460
rect 2953 456 2957 460
rect 2999 489 3003 493
rect 3005 489 3009 493
rect 3011 489 3015 493
rect 3017 489 3021 493
rect 3023 489 3027 493
rect 3029 489 3033 493
rect 3035 489 3039 493
rect 2999 471 3003 475
rect 3005 471 3009 475
rect 3011 471 3015 475
rect 3017 471 3021 475
rect 3023 471 3027 475
rect 3029 471 3033 475
rect 3035 471 3039 475
rect 2991 456 2995 460
rect 3001 456 3005 460
rect 2910 445 2914 449
rect 2916 445 2920 449
rect 2922 445 2926 449
rect 2928 445 2932 449
rect 2934 445 2938 449
rect 2910 439 2914 443
rect 2916 439 2920 443
rect 2922 439 2926 443
rect 2928 439 2932 443
rect 2934 439 2938 443
rect 2910 433 2914 437
rect 2916 433 2920 437
rect 2922 433 2926 437
rect 2928 433 2932 437
rect 2934 433 2938 437
rect 2910 427 2914 431
rect 2916 427 2920 431
rect 2922 427 2926 431
rect 2928 427 2932 431
rect 2934 427 2938 431
rect 2910 420 2914 424
rect 2916 420 2920 424
rect 2922 420 2926 424
rect 2928 420 2932 424
rect 2934 420 2938 424
rect 2910 414 2914 418
rect 2916 414 2920 418
rect 2922 414 2926 418
rect 2928 414 2932 418
rect 2934 414 2938 418
rect 3010 445 3014 449
rect 3016 445 3020 449
rect 3022 445 3026 449
rect 3028 445 3032 449
rect 3034 445 3038 449
rect 3010 439 3014 443
rect 3016 439 3020 443
rect 3022 439 3026 443
rect 3028 439 3032 443
rect 3034 439 3038 443
rect 3010 433 3014 437
rect 3016 433 3020 437
rect 3022 433 3026 437
rect 3028 433 3032 437
rect 3034 433 3038 437
rect 3010 427 3014 431
rect 3016 427 3020 431
rect 3022 427 3026 431
rect 3028 427 3032 431
rect 3034 427 3038 431
rect 3010 420 3014 424
rect 3016 420 3020 424
rect 3022 420 3026 424
rect 3028 420 3032 424
rect 3034 420 3038 424
rect 3010 414 3014 418
rect 3016 414 3020 418
rect 3022 414 3026 418
rect 3028 414 3032 418
rect 3034 414 3038 418
rect 2909 397 2913 401
rect 2915 397 2919 401
rect 2921 397 2925 401
rect 2927 397 2931 401
rect 2933 397 2937 401
rect 2939 397 2943 401
rect 2945 397 2949 401
rect 2909 384 2913 388
rect 2915 384 2919 388
rect 2921 384 2925 388
rect 2927 384 2931 388
rect 2933 384 2937 388
rect 2939 384 2943 388
rect 2945 384 2949 388
rect 2999 397 3003 401
rect 3005 397 3009 401
rect 3011 397 3015 401
rect 3017 397 3021 401
rect 3023 397 3027 401
rect 3029 397 3033 401
rect 3035 397 3039 401
rect 2999 384 3003 388
rect 3005 384 3009 388
rect 3011 384 3015 388
rect 3017 384 3021 388
rect 3023 384 3027 388
rect 3029 384 3033 388
rect 3035 384 3039 388
rect 3383 489 3387 493
rect 3389 489 3393 493
rect 3395 489 3399 493
rect 3401 489 3405 493
rect 3407 489 3411 493
rect 3413 489 3417 493
rect 3419 489 3423 493
rect 3383 471 3387 475
rect 3389 471 3393 475
rect 3395 471 3399 475
rect 3401 471 3405 475
rect 3407 471 3411 475
rect 3413 471 3417 475
rect 3419 471 3423 475
rect 3417 456 3421 460
rect 3427 456 3431 460
rect 3473 489 3477 493
rect 3479 489 3483 493
rect 3485 489 3489 493
rect 3491 489 3495 493
rect 3497 489 3501 493
rect 3503 489 3507 493
rect 3509 489 3513 493
rect 3473 471 3477 475
rect 3479 471 3483 475
rect 3485 471 3489 475
rect 3491 471 3495 475
rect 3497 471 3501 475
rect 3503 471 3507 475
rect 3509 471 3513 475
rect 3465 456 3469 460
rect 3475 456 3479 460
rect 3384 445 3388 449
rect 3390 445 3394 449
rect 3396 445 3400 449
rect 3402 445 3406 449
rect 3408 445 3412 449
rect 3384 439 3388 443
rect 3390 439 3394 443
rect 3396 439 3400 443
rect 3402 439 3406 443
rect 3408 439 3412 443
rect 3384 433 3388 437
rect 3390 433 3394 437
rect 3396 433 3400 437
rect 3402 433 3406 437
rect 3408 433 3412 437
rect 3384 427 3388 431
rect 3390 427 3394 431
rect 3396 427 3400 431
rect 3402 427 3406 431
rect 3408 427 3412 431
rect 3384 420 3388 424
rect 3390 420 3394 424
rect 3396 420 3400 424
rect 3402 420 3406 424
rect 3408 420 3412 424
rect 3384 414 3388 418
rect 3390 414 3394 418
rect 3396 414 3400 418
rect 3402 414 3406 418
rect 3408 414 3412 418
rect 3484 445 3488 449
rect 3490 445 3494 449
rect 3496 445 3500 449
rect 3502 445 3506 449
rect 3508 445 3512 449
rect 3484 439 3488 443
rect 3490 439 3494 443
rect 3496 439 3500 443
rect 3502 439 3506 443
rect 3508 439 3512 443
rect 3484 433 3488 437
rect 3490 433 3494 437
rect 3496 433 3500 437
rect 3502 433 3506 437
rect 3508 433 3512 437
rect 3484 427 3488 431
rect 3490 427 3494 431
rect 3496 427 3500 431
rect 3502 427 3506 431
rect 3508 427 3512 431
rect 3484 420 3488 424
rect 3490 420 3494 424
rect 3496 420 3500 424
rect 3502 420 3506 424
rect 3508 420 3512 424
rect 3484 414 3488 418
rect 3490 414 3494 418
rect 3496 414 3500 418
rect 3502 414 3506 418
rect 3508 414 3512 418
rect 3383 397 3387 401
rect 3389 397 3393 401
rect 3395 397 3399 401
rect 3401 397 3405 401
rect 3407 397 3411 401
rect 3413 397 3417 401
rect 3419 397 3423 401
rect 3383 384 3387 388
rect 3389 384 3393 388
rect 3395 384 3399 388
rect 3401 384 3405 388
rect 3407 384 3411 388
rect 3413 384 3417 388
rect 3419 384 3423 388
rect 3473 397 3477 401
rect 3479 397 3483 401
rect 3485 397 3489 401
rect 3491 397 3495 401
rect 3497 397 3501 401
rect 3503 397 3507 401
rect 3509 397 3513 401
rect 3473 384 3477 388
rect 3479 384 3483 388
rect 3485 384 3489 388
rect 3491 384 3495 388
rect 3497 384 3501 388
rect 3503 384 3507 388
rect 3509 384 3513 388
rect 3857 489 3861 493
rect 3863 489 3867 493
rect 3869 489 3873 493
rect 3875 489 3879 493
rect 3881 489 3885 493
rect 3887 489 3891 493
rect 3893 489 3897 493
rect 3857 471 3861 475
rect 3863 471 3867 475
rect 3869 471 3873 475
rect 3875 471 3879 475
rect 3881 471 3885 475
rect 3887 471 3891 475
rect 3893 471 3897 475
rect 3891 456 3895 460
rect 3901 456 3905 460
rect 3947 489 3951 493
rect 3953 489 3957 493
rect 3959 489 3963 493
rect 3965 489 3969 493
rect 3971 489 3975 493
rect 3977 489 3981 493
rect 3983 489 3987 493
rect 3947 471 3951 475
rect 3953 471 3957 475
rect 3959 471 3963 475
rect 3965 471 3969 475
rect 3971 471 3975 475
rect 3977 471 3981 475
rect 3983 471 3987 475
rect 3939 456 3943 460
rect 3949 456 3953 460
rect 3858 445 3862 449
rect 3864 445 3868 449
rect 3870 445 3874 449
rect 3876 445 3880 449
rect 3882 445 3886 449
rect 3858 439 3862 443
rect 3864 439 3868 443
rect 3870 439 3874 443
rect 3876 439 3880 443
rect 3882 439 3886 443
rect 3858 433 3862 437
rect 3864 433 3868 437
rect 3870 433 3874 437
rect 3876 433 3880 437
rect 3882 433 3886 437
rect 3858 427 3862 431
rect 3864 427 3868 431
rect 3870 427 3874 431
rect 3876 427 3880 431
rect 3882 427 3886 431
rect 3858 420 3862 424
rect 3864 420 3868 424
rect 3870 420 3874 424
rect 3876 420 3880 424
rect 3882 420 3886 424
rect 3858 414 3862 418
rect 3864 414 3868 418
rect 3870 414 3874 418
rect 3876 414 3880 418
rect 3882 414 3886 418
rect 3958 445 3962 449
rect 3964 445 3968 449
rect 3970 445 3974 449
rect 3976 445 3980 449
rect 3982 445 3986 449
rect 3958 439 3962 443
rect 3964 439 3968 443
rect 3970 439 3974 443
rect 3976 439 3980 443
rect 3982 439 3986 443
rect 3958 433 3962 437
rect 3964 433 3968 437
rect 3970 433 3974 437
rect 3976 433 3980 437
rect 3982 433 3986 437
rect 3958 427 3962 431
rect 3964 427 3968 431
rect 3970 427 3974 431
rect 3976 427 3980 431
rect 3982 427 3986 431
rect 3958 420 3962 424
rect 3964 420 3968 424
rect 3970 420 3974 424
rect 3976 420 3980 424
rect 3982 420 3986 424
rect 3958 414 3962 418
rect 3964 414 3968 418
rect 3970 414 3974 418
rect 3976 414 3980 418
rect 3982 414 3986 418
rect 3857 397 3861 401
rect 3863 397 3867 401
rect 3869 397 3873 401
rect 3875 397 3879 401
rect 3881 397 3885 401
rect 3887 397 3891 401
rect 3893 397 3897 401
rect 3857 384 3861 388
rect 3863 384 3867 388
rect 3869 384 3873 388
rect 3875 384 3879 388
rect 3881 384 3885 388
rect 3887 384 3891 388
rect 3893 384 3897 388
rect 3947 397 3951 401
rect 3953 397 3957 401
rect 3959 397 3963 401
rect 3965 397 3969 401
rect 3971 397 3975 401
rect 3977 397 3981 401
rect 3983 397 3987 401
rect 3947 384 3951 388
rect 3953 384 3957 388
rect 3959 384 3963 388
rect 3965 384 3969 388
rect 3971 384 3975 388
rect 3977 384 3981 388
rect 3983 384 3987 388
rect 4331 489 4335 493
rect 4337 489 4341 493
rect 4343 489 4347 493
rect 4349 489 4353 493
rect 4355 489 4359 493
rect 4361 489 4365 493
rect 4367 489 4371 493
rect 4331 471 4335 475
rect 4337 471 4341 475
rect 4343 471 4347 475
rect 4349 471 4353 475
rect 4355 471 4359 475
rect 4361 471 4365 475
rect 4367 471 4371 475
rect 4365 456 4369 460
rect 4375 456 4379 460
rect 4421 489 4425 493
rect 4427 489 4431 493
rect 4433 489 4437 493
rect 4439 489 4443 493
rect 4445 489 4449 493
rect 4451 489 4455 493
rect 4457 489 4461 493
rect 4421 471 4425 475
rect 4427 471 4431 475
rect 4433 471 4437 475
rect 4439 471 4443 475
rect 4445 471 4449 475
rect 4451 471 4455 475
rect 4457 471 4461 475
rect 4413 456 4417 460
rect 4423 456 4427 460
rect 4332 445 4336 449
rect 4338 445 4342 449
rect 4344 445 4348 449
rect 4350 445 4354 449
rect 4356 445 4360 449
rect 4332 439 4336 443
rect 4338 439 4342 443
rect 4344 439 4348 443
rect 4350 439 4354 443
rect 4356 439 4360 443
rect 4332 433 4336 437
rect 4338 433 4342 437
rect 4344 433 4348 437
rect 4350 433 4354 437
rect 4356 433 4360 437
rect 4332 427 4336 431
rect 4338 427 4342 431
rect 4344 427 4348 431
rect 4350 427 4354 431
rect 4356 427 4360 431
rect 4332 420 4336 424
rect 4338 420 4342 424
rect 4344 420 4348 424
rect 4350 420 4354 424
rect 4356 420 4360 424
rect 4332 414 4336 418
rect 4338 414 4342 418
rect 4344 414 4348 418
rect 4350 414 4354 418
rect 4356 414 4360 418
rect 4432 445 4436 449
rect 4438 445 4442 449
rect 4444 445 4448 449
rect 4450 445 4454 449
rect 4456 445 4460 449
rect 4432 439 4436 443
rect 4438 439 4442 443
rect 4444 439 4448 443
rect 4450 439 4454 443
rect 4456 439 4460 443
rect 4432 433 4436 437
rect 4438 433 4442 437
rect 4444 433 4448 437
rect 4450 433 4454 437
rect 4456 433 4460 437
rect 4432 427 4436 431
rect 4438 427 4442 431
rect 4444 427 4448 431
rect 4450 427 4454 431
rect 4456 427 4460 431
rect 4432 420 4436 424
rect 4438 420 4442 424
rect 4444 420 4448 424
rect 4450 420 4454 424
rect 4456 420 4460 424
rect 4432 414 4436 418
rect 4438 414 4442 418
rect 4444 414 4448 418
rect 4450 414 4454 418
rect 4456 414 4460 418
rect 4331 397 4335 401
rect 4337 397 4341 401
rect 4343 397 4347 401
rect 4349 397 4353 401
rect 4355 397 4359 401
rect 4361 397 4365 401
rect 4367 397 4371 401
rect 4331 384 4335 388
rect 4337 384 4341 388
rect 4343 384 4347 388
rect 4349 384 4353 388
rect 4355 384 4359 388
rect 4361 384 4365 388
rect 4367 384 4371 388
rect 4421 397 4425 401
rect 4427 397 4431 401
rect 4433 397 4437 401
rect 4439 397 4443 401
rect 4445 397 4449 401
rect 4451 397 4455 401
rect 4457 397 4461 401
rect 4421 384 4425 388
rect 4427 384 4431 388
rect 4433 384 4437 388
rect 4439 384 4443 388
rect 4445 384 4449 388
rect 4451 384 4455 388
rect 4457 384 4461 388
rect 321 249 325 253
rect 327 249 331 253
rect 333 249 337 253
rect 339 249 343 253
rect 345 249 349 253
rect 351 249 355 253
rect 321 237 325 241
rect 327 237 331 241
rect 333 237 337 241
rect 339 237 343 241
rect 345 237 349 241
rect 351 237 355 241
rect 321 225 325 229
rect 327 225 331 229
rect 333 225 337 229
rect 339 225 343 229
rect 345 225 349 229
rect 351 225 355 229
rect 4645 249 4649 253
rect 4651 249 4655 253
rect 4657 249 4661 253
rect 4663 249 4667 253
rect 4669 249 4673 253
rect 4675 249 4679 253
rect 4645 237 4649 241
rect 4651 237 4655 241
rect 4657 237 4661 241
rect 4663 237 4667 241
rect 4669 237 4673 241
rect 4675 237 4679 241
rect 4645 225 4649 229
rect 4651 225 4655 229
rect 4657 225 4661 229
rect 4663 225 4667 229
rect 4669 225 4673 229
rect 4675 225 4679 229
<< electrodecap >>
rect 465 496 668 501
rect 718 496 964 501
rect 1014 496 1142 501
rect 1192 496 1438 501
rect 1488 496 1616 501
rect 1666 496 1912 501
rect 1962 496 2090 501
rect 2140 496 2386 501
rect 2436 496 2564 501
rect 2614 496 2860 501
rect 2910 496 3038 501
rect 3088 496 3334 501
rect 3384 496 3512 501
rect 3562 496 3808 501
rect 3858 496 3986 501
rect 4036 496 4282 501
rect 4332 496 4535 501
rect 465 465 4535 496
rect 454 454 4546 462
rect 411 411 4589 451
rect 376 381 4624 408
rect 376 376 490 381
rect 540 376 668 381
rect 718 376 964 381
rect 1014 376 1142 381
rect 1192 376 1438 381
rect 1488 376 1616 381
rect 1666 376 1912 381
rect 1962 376 2090 381
rect 2140 376 2386 381
rect 2436 376 2564 381
rect 2614 376 2860 381
rect 2910 376 3038 381
rect 3088 376 3334 381
rect 3384 376 3512 381
rect 3562 376 3808 381
rect 3858 376 3986 381
rect 4036 376 4282 381
rect 4332 376 4460 381
rect 4510 376 4624 381
rect 12 353 315 358
rect 4685 353 4988 358
rect 12 318 353 353
rect 4647 318 4988 353
rect 12 315 358 318
rect 315 12 358 315
rect 4642 315 4988 318
rect 4642 12 4685 315
<< psubstratepdiff >>
rect 2 369 4998 370
rect 2 365 5 369
rect 9 365 11 369
rect 15 365 17 369
rect 21 365 23 369
rect 27 365 29 369
rect 33 365 35 369
rect 39 365 41 369
rect 45 365 47 369
rect 51 365 53 369
rect 57 365 59 369
rect 63 365 65 369
rect 69 365 71 369
rect 75 365 77 369
rect 81 365 83 369
rect 87 365 89 369
rect 93 365 95 369
rect 99 365 101 369
rect 105 365 107 369
rect 111 365 113 369
rect 117 365 119 369
rect 123 365 125 369
rect 129 365 131 369
rect 135 365 137 369
rect 141 365 143 369
rect 147 365 149 369
rect 153 365 155 369
rect 159 365 161 369
rect 165 365 167 369
rect 171 365 173 369
rect 177 365 179 369
rect 183 365 185 369
rect 189 365 191 369
rect 195 365 197 369
rect 201 365 203 369
rect 207 365 209 369
rect 213 365 215 369
rect 219 365 221 369
rect 225 365 227 369
rect 231 365 233 369
rect 237 365 239 369
rect 243 365 245 369
rect 249 365 251 369
rect 255 365 257 369
rect 261 365 263 369
rect 267 365 269 369
rect 273 365 275 369
rect 279 365 281 369
rect 285 365 287 369
rect 291 365 293 369
rect 297 365 299 369
rect 303 365 305 369
rect 309 365 311 369
rect 315 365 317 369
rect 321 365 323 369
rect 327 365 329 369
rect 333 365 335 369
rect 339 365 341 369
rect 345 365 347 369
rect 351 365 353 369
rect 357 365 359 369
rect 363 365 365 369
rect 369 365 371 369
rect 375 365 377 369
rect 381 365 383 369
rect 387 365 389 369
rect 393 365 395 369
rect 399 365 401 369
rect 405 365 407 369
rect 411 365 413 369
rect 417 365 419 369
rect 423 365 425 369
rect 429 365 431 369
rect 435 365 437 369
rect 441 365 443 369
rect 447 365 449 369
rect 453 365 455 369
rect 459 365 461 369
rect 465 365 467 369
rect 471 365 473 369
rect 477 365 479 369
rect 483 365 485 369
rect 489 365 491 369
rect 495 365 497 369
rect 501 365 503 369
rect 507 365 509 369
rect 513 365 515 369
rect 519 365 521 369
rect 525 365 527 369
rect 531 365 533 369
rect 537 365 539 369
rect 543 365 545 369
rect 549 365 551 369
rect 555 365 557 369
rect 561 365 563 369
rect 567 365 569 369
rect 573 365 575 369
rect 579 365 581 369
rect 585 365 587 369
rect 591 365 617 369
rect 621 365 623 369
rect 627 365 629 369
rect 633 365 635 369
rect 639 365 641 369
rect 645 365 647 369
rect 651 365 653 369
rect 657 365 659 369
rect 663 365 665 369
rect 669 365 671 369
rect 675 365 677 369
rect 681 365 683 369
rect 687 365 689 369
rect 693 365 695 369
rect 699 365 701 369
rect 705 365 707 369
rect 711 365 713 369
rect 717 365 719 369
rect 723 365 725 369
rect 729 365 731 369
rect 735 365 737 369
rect 741 365 743 369
rect 747 365 749 369
rect 753 365 755 369
rect 759 365 761 369
rect 765 365 767 369
rect 771 365 773 369
rect 777 365 779 369
rect 783 365 785 369
rect 789 365 791 369
rect 795 365 797 369
rect 801 365 803 369
rect 807 365 809 369
rect 813 365 815 369
rect 819 365 821 369
rect 825 365 827 369
rect 831 365 833 369
rect 837 365 839 369
rect 843 365 845 369
rect 849 365 851 369
rect 855 365 857 369
rect 861 365 863 369
rect 867 365 869 369
rect 873 365 875 369
rect 879 365 881 369
rect 885 365 887 369
rect 891 365 893 369
rect 897 365 899 369
rect 903 365 905 369
rect 909 365 911 369
rect 915 365 917 369
rect 921 365 923 369
rect 927 365 929 369
rect 933 365 935 369
rect 939 365 941 369
rect 945 365 947 369
rect 951 365 953 369
rect 957 365 959 369
rect 963 365 965 369
rect 969 365 971 369
rect 975 365 977 369
rect 981 365 983 369
rect 987 365 989 369
rect 993 365 995 369
rect 999 365 1001 369
rect 1005 365 1007 369
rect 1011 365 1013 369
rect 1017 365 1019 369
rect 1023 365 1025 369
rect 1029 365 1031 369
rect 1035 365 1037 369
rect 1041 365 1043 369
rect 1047 365 1049 369
rect 1053 365 1055 369
rect 1059 365 1061 369
rect 1065 365 1091 369
rect 1095 365 1097 369
rect 1101 365 1103 369
rect 1107 365 1109 369
rect 1113 365 1115 369
rect 1119 365 1121 369
rect 1125 365 1127 369
rect 1131 365 1133 369
rect 1137 365 1139 369
rect 1143 365 1145 369
rect 1149 365 1151 369
rect 1155 365 1157 369
rect 1161 365 1163 369
rect 1167 365 1169 369
rect 1173 365 1175 369
rect 1179 365 1181 369
rect 1185 365 1187 369
rect 1191 365 1193 369
rect 1197 365 1199 369
rect 1203 365 1205 369
rect 1209 365 1211 369
rect 1215 365 1217 369
rect 1221 365 1223 369
rect 1227 365 1229 369
rect 1233 365 1235 369
rect 1239 365 1241 369
rect 1245 365 1247 369
rect 1251 365 1253 369
rect 1257 365 1259 369
rect 1263 365 1265 369
rect 1269 365 1271 369
rect 1275 365 1277 369
rect 1281 365 1283 369
rect 1287 365 1289 369
rect 1293 365 1295 369
rect 1299 365 1301 369
rect 1305 365 1307 369
rect 1311 365 1313 369
rect 1317 365 1319 369
rect 1323 365 1325 369
rect 1329 365 1331 369
rect 1335 365 1337 369
rect 1341 365 1343 369
rect 1347 365 1349 369
rect 1353 365 1355 369
rect 1359 365 1361 369
rect 1365 365 1367 369
rect 1371 365 1373 369
rect 1377 365 1379 369
rect 1383 365 1385 369
rect 1389 365 1391 369
rect 1395 365 1397 369
rect 1401 365 1403 369
rect 1407 365 1409 369
rect 1413 365 1415 369
rect 1419 365 1421 369
rect 1425 365 1427 369
rect 1431 365 1433 369
rect 1437 365 1439 369
rect 1443 365 1445 369
rect 1449 365 1451 369
rect 1455 365 1457 369
rect 1461 365 1463 369
rect 1467 365 1469 369
rect 1473 365 1475 369
rect 1479 365 1481 369
rect 1485 365 1487 369
rect 1491 365 1493 369
rect 1497 365 1499 369
rect 1503 365 1505 369
rect 1509 365 1511 369
rect 1515 365 1517 369
rect 1521 365 1523 369
rect 1527 365 1529 369
rect 1533 365 1535 369
rect 1539 365 1565 369
rect 1569 365 1571 369
rect 1575 365 1577 369
rect 1581 365 1583 369
rect 1587 365 1589 369
rect 1593 365 1595 369
rect 1599 365 1601 369
rect 1605 365 1607 369
rect 1611 365 1613 369
rect 1617 365 1619 369
rect 1623 365 1625 369
rect 1629 365 1631 369
rect 1635 365 1637 369
rect 1641 365 1643 369
rect 1647 365 1649 369
rect 1653 365 1655 369
rect 1659 365 1661 369
rect 1665 365 1667 369
rect 1671 365 1673 369
rect 1677 365 1679 369
rect 1683 365 1685 369
rect 1689 365 1691 369
rect 1695 365 1697 369
rect 1701 365 1703 369
rect 1707 365 1709 369
rect 1713 365 1715 369
rect 1719 365 1721 369
rect 1725 365 1727 369
rect 1731 365 1733 369
rect 1737 365 1739 369
rect 1743 365 1745 369
rect 1749 365 1751 369
rect 1755 365 1757 369
rect 1761 365 1763 369
rect 1767 365 1769 369
rect 1773 365 1775 369
rect 1779 365 1781 369
rect 1785 365 1787 369
rect 1791 365 1793 369
rect 1797 365 1799 369
rect 1803 365 1805 369
rect 1809 365 1811 369
rect 1815 365 1817 369
rect 1821 365 1823 369
rect 1827 365 1829 369
rect 1833 365 1835 369
rect 1839 365 1841 369
rect 1845 365 1847 369
rect 1851 365 1853 369
rect 1857 365 1859 369
rect 1863 365 1865 369
rect 1869 365 1871 369
rect 1875 365 1877 369
rect 1881 365 1883 369
rect 1887 365 1889 369
rect 1893 365 1895 369
rect 1899 365 1901 369
rect 1905 365 1907 369
rect 1911 365 1913 369
rect 1917 365 1919 369
rect 1923 365 1925 369
rect 1929 365 1931 369
rect 1935 365 1937 369
rect 1941 365 1943 369
rect 1947 365 1949 369
rect 1953 365 1955 369
rect 1959 365 1961 369
rect 1965 365 1967 369
rect 1971 365 1973 369
rect 1977 365 1979 369
rect 1983 365 1985 369
rect 1989 365 1991 369
rect 1995 365 1997 369
rect 2001 365 2003 369
rect 2007 365 2009 369
rect 2013 365 2039 369
rect 2043 365 2045 369
rect 2049 365 2051 369
rect 2055 365 2057 369
rect 2061 365 2063 369
rect 2067 365 2069 369
rect 2073 365 2075 369
rect 2079 365 2081 369
rect 2085 365 2087 369
rect 2091 365 2093 369
rect 2097 365 2099 369
rect 2103 365 2105 369
rect 2109 365 2111 369
rect 2115 365 2117 369
rect 2121 365 2123 369
rect 2127 365 2129 369
rect 2133 365 2135 369
rect 2139 365 2141 369
rect 2145 365 2147 369
rect 2151 365 2153 369
rect 2157 365 2159 369
rect 2163 365 2165 369
rect 2169 365 2171 369
rect 2175 365 2177 369
rect 2181 365 2183 369
rect 2187 365 2189 369
rect 2193 365 2195 369
rect 2199 365 2201 369
rect 2205 365 2207 369
rect 2211 365 2213 369
rect 2217 365 2219 369
rect 2223 365 2225 369
rect 2229 365 2231 369
rect 2235 365 2237 369
rect 2241 365 2243 369
rect 2247 365 2249 369
rect 2253 365 2255 369
rect 2259 365 2261 369
rect 2265 365 2267 369
rect 2271 365 2273 369
rect 2277 365 2279 369
rect 2283 365 2285 369
rect 2289 365 2291 369
rect 2295 365 2297 369
rect 2301 365 2303 369
rect 2307 365 2309 369
rect 2313 365 2315 369
rect 2319 365 2321 369
rect 2325 365 2327 369
rect 2331 365 2333 369
rect 2337 365 2339 369
rect 2343 365 2345 369
rect 2349 365 2351 369
rect 2355 365 2357 369
rect 2361 365 2363 369
rect 2367 365 2369 369
rect 2373 365 2375 369
rect 2379 365 2381 369
rect 2385 365 2387 369
rect 2391 365 2393 369
rect 2397 365 2399 369
rect 2403 365 2405 369
rect 2409 365 2411 369
rect 2415 365 2417 369
rect 2421 365 2423 369
rect 2427 365 2429 369
rect 2433 365 2435 369
rect 2439 365 2441 369
rect 2445 365 2447 369
rect 2451 365 2453 369
rect 2457 365 2459 369
rect 2463 365 2465 369
rect 2469 365 2471 369
rect 2475 365 2477 369
rect 2481 365 2483 369
rect 2487 365 2513 369
rect 2517 365 2519 369
rect 2523 365 2525 369
rect 2529 365 2531 369
rect 2535 365 2537 369
rect 2541 365 2543 369
rect 2547 365 2549 369
rect 2553 365 2555 369
rect 2559 365 2561 369
rect 2565 365 2567 369
rect 2571 365 2573 369
rect 2577 365 2579 369
rect 2583 365 2585 369
rect 2589 365 2591 369
rect 2595 365 2597 369
rect 2601 365 2603 369
rect 2607 365 2609 369
rect 2613 365 2615 369
rect 2619 365 2621 369
rect 2625 365 2627 369
rect 2631 365 2633 369
rect 2637 365 2639 369
rect 2643 365 2645 369
rect 2649 365 2651 369
rect 2655 365 2657 369
rect 2661 365 2663 369
rect 2667 365 2669 369
rect 2673 365 2675 369
rect 2679 365 2681 369
rect 2685 365 2687 369
rect 2691 365 2693 369
rect 2697 365 2699 369
rect 2703 365 2705 369
rect 2709 365 2711 369
rect 2715 365 2717 369
rect 2721 365 2723 369
rect 2727 365 2729 369
rect 2733 365 2735 369
rect 2739 365 2741 369
rect 2745 365 2747 369
rect 2751 365 2753 369
rect 2757 365 2759 369
rect 2763 365 2765 369
rect 2769 365 2771 369
rect 2775 365 2777 369
rect 2781 365 2783 369
rect 2787 365 2789 369
rect 2793 365 2795 369
rect 2799 365 2801 369
rect 2805 365 2807 369
rect 2811 365 2813 369
rect 2817 365 2819 369
rect 2823 365 2825 369
rect 2829 365 2831 369
rect 2835 365 2837 369
rect 2841 365 2843 369
rect 2847 365 2849 369
rect 2853 365 2855 369
rect 2859 365 2861 369
rect 2865 365 2867 369
rect 2871 365 2873 369
rect 2877 365 2879 369
rect 2883 365 2885 369
rect 2889 365 2891 369
rect 2895 365 2897 369
rect 2901 365 2903 369
rect 2907 365 2909 369
rect 2913 365 2915 369
rect 2919 365 2921 369
rect 2925 365 2927 369
rect 2931 365 2933 369
rect 2937 365 2939 369
rect 2943 365 2945 369
rect 2949 365 2951 369
rect 2955 365 2957 369
rect 2961 365 2987 369
rect 2991 365 2993 369
rect 2997 365 2999 369
rect 3003 365 3005 369
rect 3009 365 3011 369
rect 3015 365 3017 369
rect 3021 365 3023 369
rect 3027 365 3029 369
rect 3033 365 3035 369
rect 3039 365 3041 369
rect 3045 365 3047 369
rect 3051 365 3053 369
rect 3057 365 3059 369
rect 3063 365 3065 369
rect 3069 365 3071 369
rect 3075 365 3077 369
rect 3081 365 3083 369
rect 3087 365 3089 369
rect 3093 365 3095 369
rect 3099 365 3101 369
rect 3105 365 3107 369
rect 3111 365 3113 369
rect 3117 365 3119 369
rect 3123 365 3125 369
rect 3129 365 3131 369
rect 3135 365 3137 369
rect 3141 365 3143 369
rect 3147 365 3149 369
rect 3153 365 3155 369
rect 3159 365 3161 369
rect 3165 365 3167 369
rect 3171 365 3173 369
rect 3177 365 3179 369
rect 3183 365 3185 369
rect 3189 365 3191 369
rect 3195 365 3197 369
rect 3201 365 3203 369
rect 3207 365 3209 369
rect 3213 365 3215 369
rect 3219 365 3221 369
rect 3225 365 3227 369
rect 3231 365 3233 369
rect 3237 365 3239 369
rect 3243 365 3245 369
rect 3249 365 3251 369
rect 3255 365 3257 369
rect 3261 365 3263 369
rect 3267 365 3269 369
rect 3273 365 3275 369
rect 3279 365 3281 369
rect 3285 365 3287 369
rect 3291 365 3293 369
rect 3297 365 3299 369
rect 3303 365 3305 369
rect 3309 365 3311 369
rect 3315 365 3317 369
rect 3321 365 3323 369
rect 3327 365 3329 369
rect 3333 365 3335 369
rect 3339 365 3341 369
rect 3345 365 3347 369
rect 3351 365 3353 369
rect 3357 365 3359 369
rect 3363 365 3365 369
rect 3369 365 3371 369
rect 3375 365 3377 369
rect 3381 365 3383 369
rect 3387 365 3389 369
rect 3393 365 3395 369
rect 3399 365 3401 369
rect 3405 365 3407 369
rect 3411 365 3413 369
rect 3417 365 3419 369
rect 3423 365 3425 369
rect 3429 365 3431 369
rect 3435 365 3461 369
rect 3465 365 3467 369
rect 3471 365 3473 369
rect 3477 365 3479 369
rect 3483 365 3485 369
rect 3489 365 3491 369
rect 3495 365 3497 369
rect 3501 365 3503 369
rect 3507 365 3509 369
rect 3513 365 3515 369
rect 3519 365 3521 369
rect 3525 365 3527 369
rect 3531 365 3533 369
rect 3537 365 3539 369
rect 3543 365 3545 369
rect 3549 365 3551 369
rect 3555 365 3557 369
rect 3561 365 3563 369
rect 3567 365 3569 369
rect 3573 365 3575 369
rect 3579 365 3581 369
rect 3585 365 3587 369
rect 3591 365 3593 369
rect 3597 365 3599 369
rect 3603 365 3605 369
rect 3609 365 3611 369
rect 3615 365 3617 369
rect 3621 365 3623 369
rect 3627 365 3629 369
rect 3633 365 3635 369
rect 3639 365 3641 369
rect 3645 365 3647 369
rect 3651 365 3653 369
rect 3657 365 3659 369
rect 3663 365 3665 369
rect 3669 365 3671 369
rect 3675 365 3677 369
rect 3681 365 3683 369
rect 3687 365 3689 369
rect 3693 365 3695 369
rect 3699 365 3701 369
rect 3705 365 3707 369
rect 3711 365 3713 369
rect 3717 365 3719 369
rect 3723 365 3725 369
rect 3729 365 3731 369
rect 3735 365 3737 369
rect 3741 365 3743 369
rect 3747 365 3749 369
rect 3753 365 3755 369
rect 3759 365 3761 369
rect 3765 365 3767 369
rect 3771 365 3773 369
rect 3777 365 3779 369
rect 3783 365 3785 369
rect 3789 365 3791 369
rect 3795 365 3797 369
rect 3801 365 3803 369
rect 3807 365 3809 369
rect 3813 365 3815 369
rect 3819 365 3821 369
rect 3825 365 3827 369
rect 3831 365 3833 369
rect 3837 365 3839 369
rect 3843 365 3845 369
rect 3849 365 3851 369
rect 3855 365 3857 369
rect 3861 365 3863 369
rect 3867 365 3869 369
rect 3873 365 3875 369
rect 3879 365 3881 369
rect 3885 365 3887 369
rect 3891 365 3893 369
rect 3897 365 3899 369
rect 3903 365 3905 369
rect 3909 365 3935 369
rect 3939 365 3941 369
rect 3945 365 3947 369
rect 3951 365 3953 369
rect 3957 365 3959 369
rect 3963 365 3965 369
rect 3969 365 3971 369
rect 3975 365 3977 369
rect 3981 365 3983 369
rect 3987 365 3989 369
rect 3993 365 3995 369
rect 3999 365 4001 369
rect 4005 365 4007 369
rect 4011 365 4013 369
rect 4017 365 4019 369
rect 4023 365 4025 369
rect 4029 365 4031 369
rect 4035 365 4037 369
rect 4041 365 4043 369
rect 4047 365 4049 369
rect 4053 365 4055 369
rect 4059 365 4061 369
rect 4065 365 4067 369
rect 4071 365 4073 369
rect 4077 365 4079 369
rect 4083 365 4085 369
rect 4089 365 4091 369
rect 4095 365 4097 369
rect 4101 365 4103 369
rect 4107 365 4109 369
rect 4113 365 4115 369
rect 4119 365 4121 369
rect 4125 365 4127 369
rect 4131 365 4133 369
rect 4137 365 4139 369
rect 4143 365 4145 369
rect 4149 365 4151 369
rect 4155 365 4157 369
rect 4161 365 4163 369
rect 4167 365 4169 369
rect 4173 365 4175 369
rect 4179 365 4181 369
rect 4185 365 4187 369
rect 4191 365 4193 369
rect 4197 365 4199 369
rect 4203 365 4205 369
rect 4209 365 4211 369
rect 4215 365 4217 369
rect 4221 365 4223 369
rect 4227 365 4229 369
rect 4233 365 4235 369
rect 4239 365 4241 369
rect 4245 365 4247 369
rect 4251 365 4253 369
rect 4257 365 4259 369
rect 4263 365 4265 369
rect 4269 365 4271 369
rect 4275 365 4277 369
rect 4281 365 4283 369
rect 4287 365 4289 369
rect 4293 365 4295 369
rect 4299 365 4301 369
rect 4305 365 4307 369
rect 4311 365 4313 369
rect 4317 365 4319 369
rect 4323 365 4325 369
rect 4329 365 4331 369
rect 4335 365 4337 369
rect 4341 365 4343 369
rect 4347 365 4349 369
rect 4353 365 4355 369
rect 4359 365 4361 369
rect 4365 365 4367 369
rect 4371 365 4373 369
rect 4377 365 4379 369
rect 4383 365 4409 369
rect 4413 365 4415 369
rect 4419 365 4421 369
rect 4425 365 4427 369
rect 4431 365 4433 369
rect 4437 365 4439 369
rect 4443 365 4445 369
rect 4449 365 4451 369
rect 4455 365 4457 369
rect 4461 365 4463 369
rect 4467 365 4469 369
rect 4473 365 4475 369
rect 4479 365 4481 369
rect 4485 365 4487 369
rect 4491 365 4493 369
rect 4497 365 4499 369
rect 4503 365 4505 369
rect 4509 365 4511 369
rect 4515 365 4517 369
rect 4521 365 4523 369
rect 4527 365 4529 369
rect 4533 365 4535 369
rect 4539 365 4541 369
rect 4545 365 4547 369
rect 4551 365 4553 369
rect 4557 365 4559 369
rect 4563 365 4565 369
rect 4569 365 4571 369
rect 4575 365 4577 369
rect 4581 365 4583 369
rect 4587 365 4589 369
rect 4593 365 4595 369
rect 4599 365 4601 369
rect 4605 365 4607 369
rect 4611 365 4613 369
rect 4617 365 4619 369
rect 4623 365 4625 369
rect 4629 365 4631 369
rect 4635 365 4637 369
rect 4641 365 4643 369
rect 4647 365 4649 369
rect 4653 365 4655 369
rect 4659 365 4661 369
rect 4665 365 4667 369
rect 4671 365 4673 369
rect 4677 365 4679 369
rect 4683 365 4685 369
rect 4689 365 4691 369
rect 4695 365 4697 369
rect 4701 365 4703 369
rect 4707 365 4709 369
rect 4713 365 4715 369
rect 4719 365 4721 369
rect 4725 365 4727 369
rect 4731 365 4733 369
rect 4737 365 4739 369
rect 4743 365 4745 369
rect 4749 365 4751 369
rect 4755 365 4757 369
rect 4761 365 4763 369
rect 4767 365 4769 369
rect 4773 365 4775 369
rect 4779 365 4781 369
rect 4785 365 4787 369
rect 4791 365 4793 369
rect 4797 365 4799 369
rect 4803 365 4805 369
rect 4809 365 4811 369
rect 4815 365 4817 369
rect 4821 365 4823 369
rect 4827 365 4829 369
rect 4833 365 4835 369
rect 4839 365 4841 369
rect 4845 365 4847 369
rect 4851 365 4853 369
rect 4857 365 4859 369
rect 4863 365 4865 369
rect 4869 365 4871 369
rect 4875 365 4877 369
rect 4881 365 4883 369
rect 4887 365 4889 369
rect 4893 365 4895 369
rect 4899 365 4901 369
rect 4905 365 4907 369
rect 4911 365 4913 369
rect 4917 365 4919 369
rect 4923 365 4925 369
rect 4929 365 4931 369
rect 4935 365 4937 369
rect 4941 365 4943 369
rect 4947 365 4949 369
rect 4953 365 4955 369
rect 4959 365 4961 369
rect 4965 365 4967 369
rect 4971 365 4973 369
rect 4977 365 4979 369
rect 4983 365 4985 369
rect 4989 365 4991 369
rect 4995 365 4998 369
rect 2 364 4998 365
rect 364 363 370 364
rect 364 359 365 363
rect 369 359 370 363
rect 364 357 370 359
rect 364 353 365 357
rect 369 353 370 357
rect 364 351 370 353
rect 364 347 365 351
rect 369 347 370 351
rect 364 345 370 347
rect 364 341 365 345
rect 369 341 370 345
rect 364 339 370 341
rect 364 335 365 339
rect 369 335 370 339
rect 364 333 370 335
rect 364 329 365 333
rect 369 329 370 333
rect 364 327 370 329
rect 364 323 365 327
rect 369 323 370 327
rect 364 321 370 323
rect 364 317 365 321
rect 369 317 370 321
rect 364 315 370 317
rect 364 311 365 315
rect 369 311 370 315
rect 364 309 370 311
rect 364 305 365 309
rect 369 305 370 309
rect 364 303 370 305
rect 364 299 365 303
rect 369 299 370 303
rect 364 297 370 299
rect 364 293 365 297
rect 369 293 370 297
rect 364 291 370 293
rect 364 287 365 291
rect 369 287 370 291
rect 364 285 370 287
rect 364 281 365 285
rect 369 281 370 285
rect 364 279 370 281
rect 364 275 365 279
rect 369 275 370 279
rect 364 273 370 275
rect 364 269 365 273
rect 369 269 370 273
rect 364 267 370 269
rect 364 263 365 267
rect 369 263 370 267
rect 364 261 370 263
rect 364 257 365 261
rect 369 257 370 261
rect 364 255 370 257
rect 364 251 365 255
rect 369 251 370 255
rect 364 249 370 251
rect 364 245 365 249
rect 369 245 370 249
rect 364 243 370 245
rect 364 239 365 243
rect 369 239 370 243
rect 364 237 370 239
rect 364 233 365 237
rect 369 233 370 237
rect 364 231 370 233
rect 364 227 365 231
rect 369 227 370 231
rect 364 225 370 227
rect 364 221 365 225
rect 369 221 370 225
rect 364 219 370 221
rect 364 215 365 219
rect 369 215 370 219
rect 364 213 370 215
rect 364 209 365 213
rect 369 209 370 213
rect 364 207 370 209
rect 364 203 365 207
rect 369 203 370 207
rect 364 201 370 203
rect 364 197 365 201
rect 369 197 370 201
rect 364 195 370 197
rect 364 191 365 195
rect 369 191 370 195
rect 364 189 370 191
rect 364 185 365 189
rect 369 185 370 189
rect 364 183 370 185
rect 364 179 365 183
rect 369 179 370 183
rect 364 177 370 179
rect 364 173 365 177
rect 369 173 370 177
rect 364 171 370 173
rect 364 167 365 171
rect 369 167 370 171
rect 364 165 370 167
rect 364 161 365 165
rect 369 161 370 165
rect 364 159 370 161
rect 364 155 365 159
rect 369 155 370 159
rect 364 153 370 155
rect 364 149 365 153
rect 369 149 370 153
rect 364 147 370 149
rect 364 143 365 147
rect 369 143 370 147
rect 364 141 370 143
rect 364 137 365 141
rect 369 137 370 141
rect 364 135 370 137
rect 364 131 365 135
rect 369 131 370 135
rect 364 129 370 131
rect 364 125 365 129
rect 369 125 370 129
rect 364 123 370 125
rect 364 119 365 123
rect 369 119 370 123
rect 364 117 370 119
rect 364 113 365 117
rect 369 113 370 117
rect 364 111 370 113
rect 364 107 365 111
rect 369 107 370 111
rect 364 105 370 107
rect 364 101 365 105
rect 369 101 370 105
rect 364 99 370 101
rect 364 95 365 99
rect 369 95 370 99
rect 364 93 370 95
rect 364 89 365 93
rect 369 89 370 93
rect 364 87 370 89
rect 364 83 365 87
rect 369 83 370 87
rect 364 81 370 83
rect 364 77 365 81
rect 369 77 370 81
rect 364 75 370 77
rect 364 71 365 75
rect 369 71 370 75
rect 364 69 370 71
rect 364 65 365 69
rect 369 65 370 69
rect 364 63 370 65
rect 364 59 365 63
rect 369 59 370 63
rect 364 57 370 59
rect 364 53 365 57
rect 369 53 370 57
rect 364 51 370 53
rect 364 47 365 51
rect 369 47 370 51
rect 364 45 370 47
rect 364 41 365 45
rect 369 41 370 45
rect 364 39 370 41
rect 364 35 365 39
rect 369 35 370 39
rect 364 33 370 35
rect 364 29 365 33
rect 369 29 370 33
rect 364 27 370 29
rect 364 23 365 27
rect 369 23 370 27
rect 364 21 370 23
rect 364 17 365 21
rect 369 17 370 21
rect 364 15 370 17
rect 364 11 365 15
rect 369 11 370 15
rect 364 9 370 11
rect 364 5 365 9
rect 369 5 370 9
rect 364 2 370 5
rect 838 363 844 364
rect 838 359 839 363
rect 843 359 844 363
rect 838 357 844 359
rect 838 353 839 357
rect 843 353 844 357
rect 838 351 844 353
rect 838 347 839 351
rect 843 347 844 351
rect 838 345 844 347
rect 838 341 839 345
rect 843 341 844 345
rect 838 339 844 341
rect 838 335 839 339
rect 843 335 844 339
rect 838 333 844 335
rect 838 329 839 333
rect 843 329 844 333
rect 838 327 844 329
rect 838 323 839 327
rect 843 323 844 327
rect 838 321 844 323
rect 838 317 839 321
rect 843 317 844 321
rect 838 315 844 317
rect 838 311 839 315
rect 843 311 844 315
rect 838 309 844 311
rect 838 305 839 309
rect 843 305 844 309
rect 838 303 844 305
rect 838 299 839 303
rect 843 299 844 303
rect 838 297 844 299
rect 838 293 839 297
rect 843 293 844 297
rect 838 291 844 293
rect 838 287 839 291
rect 843 287 844 291
rect 838 285 844 287
rect 838 281 839 285
rect 843 281 844 285
rect 838 279 844 281
rect 838 275 839 279
rect 843 275 844 279
rect 838 273 844 275
rect 838 269 839 273
rect 843 269 844 273
rect 838 267 844 269
rect 838 263 839 267
rect 843 263 844 267
rect 838 261 844 263
rect 838 257 839 261
rect 843 257 844 261
rect 838 255 844 257
rect 838 251 839 255
rect 843 251 844 255
rect 838 249 844 251
rect 838 245 839 249
rect 843 245 844 249
rect 838 243 844 245
rect 838 239 839 243
rect 843 239 844 243
rect 838 237 844 239
rect 838 233 839 237
rect 843 233 844 237
rect 838 231 844 233
rect 838 227 839 231
rect 843 227 844 231
rect 838 225 844 227
rect 838 221 839 225
rect 843 221 844 225
rect 838 219 844 221
rect 838 215 839 219
rect 843 215 844 219
rect 838 213 844 215
rect 838 209 839 213
rect 843 209 844 213
rect 838 207 844 209
rect 838 203 839 207
rect 843 203 844 207
rect 838 201 844 203
rect 838 197 839 201
rect 843 197 844 201
rect 838 195 844 197
rect 838 191 839 195
rect 843 191 844 195
rect 838 189 844 191
rect 838 185 839 189
rect 843 185 844 189
rect 838 183 844 185
rect 838 179 839 183
rect 843 179 844 183
rect 838 177 844 179
rect 838 173 839 177
rect 843 173 844 177
rect 838 171 844 173
rect 838 167 839 171
rect 843 167 844 171
rect 838 165 844 167
rect 838 161 839 165
rect 843 161 844 165
rect 838 159 844 161
rect 838 155 839 159
rect 843 155 844 159
rect 838 153 844 155
rect 838 149 839 153
rect 843 149 844 153
rect 838 147 844 149
rect 838 143 839 147
rect 843 143 844 147
rect 838 141 844 143
rect 838 137 839 141
rect 843 137 844 141
rect 838 135 844 137
rect 838 131 839 135
rect 843 131 844 135
rect 838 129 844 131
rect 838 125 839 129
rect 843 125 844 129
rect 838 123 844 125
rect 838 119 839 123
rect 843 119 844 123
rect 838 117 844 119
rect 838 113 839 117
rect 843 113 844 117
rect 838 111 844 113
rect 838 107 839 111
rect 843 107 844 111
rect 838 105 844 107
rect 838 101 839 105
rect 843 101 844 105
rect 838 99 844 101
rect 838 95 839 99
rect 843 95 844 99
rect 838 93 844 95
rect 838 89 839 93
rect 843 89 844 93
rect 838 87 844 89
rect 838 83 839 87
rect 843 83 844 87
rect 838 81 844 83
rect 838 77 839 81
rect 843 77 844 81
rect 838 75 844 77
rect 838 71 839 75
rect 843 71 844 75
rect 838 69 844 71
rect 838 65 839 69
rect 843 65 844 69
rect 838 63 844 65
rect 838 59 839 63
rect 843 59 844 63
rect 838 57 844 59
rect 838 53 839 57
rect 843 53 844 57
rect 838 51 844 53
rect 838 47 839 51
rect 843 47 844 51
rect 838 45 844 47
rect 838 41 839 45
rect 843 41 844 45
rect 838 39 844 41
rect 838 35 839 39
rect 843 35 844 39
rect 838 33 844 35
rect 838 29 839 33
rect 843 29 844 33
rect 838 27 844 29
rect 838 23 839 27
rect 843 23 844 27
rect 838 21 844 23
rect 838 17 839 21
rect 843 17 844 21
rect 838 15 844 17
rect 838 11 839 15
rect 843 11 844 15
rect 838 9 844 11
rect 838 5 839 9
rect 843 5 844 9
rect 838 2 844 5
rect 1312 363 1318 364
rect 1312 359 1313 363
rect 1317 359 1318 363
rect 1312 357 1318 359
rect 1312 353 1313 357
rect 1317 353 1318 357
rect 1312 351 1318 353
rect 1312 347 1313 351
rect 1317 347 1318 351
rect 1312 345 1318 347
rect 1312 341 1313 345
rect 1317 341 1318 345
rect 1312 339 1318 341
rect 1312 335 1313 339
rect 1317 335 1318 339
rect 1312 333 1318 335
rect 1312 329 1313 333
rect 1317 329 1318 333
rect 1312 327 1318 329
rect 1312 323 1313 327
rect 1317 323 1318 327
rect 1312 321 1318 323
rect 1312 317 1313 321
rect 1317 317 1318 321
rect 1312 315 1318 317
rect 1312 311 1313 315
rect 1317 311 1318 315
rect 1312 309 1318 311
rect 1312 305 1313 309
rect 1317 305 1318 309
rect 1312 303 1318 305
rect 1312 299 1313 303
rect 1317 299 1318 303
rect 1312 297 1318 299
rect 1312 293 1313 297
rect 1317 293 1318 297
rect 1312 291 1318 293
rect 1312 287 1313 291
rect 1317 287 1318 291
rect 1312 285 1318 287
rect 1312 281 1313 285
rect 1317 281 1318 285
rect 1312 279 1318 281
rect 1312 275 1313 279
rect 1317 275 1318 279
rect 1312 273 1318 275
rect 1312 269 1313 273
rect 1317 269 1318 273
rect 1312 267 1318 269
rect 1312 263 1313 267
rect 1317 263 1318 267
rect 1312 261 1318 263
rect 1312 257 1313 261
rect 1317 257 1318 261
rect 1312 255 1318 257
rect 1312 251 1313 255
rect 1317 251 1318 255
rect 1312 249 1318 251
rect 1312 245 1313 249
rect 1317 245 1318 249
rect 1312 243 1318 245
rect 1312 239 1313 243
rect 1317 239 1318 243
rect 1312 237 1318 239
rect 1312 233 1313 237
rect 1317 233 1318 237
rect 1312 231 1318 233
rect 1312 227 1313 231
rect 1317 227 1318 231
rect 1312 225 1318 227
rect 1312 221 1313 225
rect 1317 221 1318 225
rect 1312 219 1318 221
rect 1312 215 1313 219
rect 1317 215 1318 219
rect 1312 213 1318 215
rect 1312 209 1313 213
rect 1317 209 1318 213
rect 1312 207 1318 209
rect 1312 203 1313 207
rect 1317 203 1318 207
rect 1312 201 1318 203
rect 1312 197 1313 201
rect 1317 197 1318 201
rect 1312 195 1318 197
rect 1312 191 1313 195
rect 1317 191 1318 195
rect 1312 189 1318 191
rect 1312 185 1313 189
rect 1317 185 1318 189
rect 1312 183 1318 185
rect 1312 179 1313 183
rect 1317 179 1318 183
rect 1312 177 1318 179
rect 1312 173 1313 177
rect 1317 173 1318 177
rect 1312 171 1318 173
rect 1312 167 1313 171
rect 1317 167 1318 171
rect 1312 165 1318 167
rect 1312 161 1313 165
rect 1317 161 1318 165
rect 1312 159 1318 161
rect 1312 155 1313 159
rect 1317 155 1318 159
rect 1312 153 1318 155
rect 1312 149 1313 153
rect 1317 149 1318 153
rect 1312 147 1318 149
rect 1312 143 1313 147
rect 1317 143 1318 147
rect 1312 141 1318 143
rect 1312 137 1313 141
rect 1317 137 1318 141
rect 1312 135 1318 137
rect 1312 131 1313 135
rect 1317 131 1318 135
rect 1312 129 1318 131
rect 1312 125 1313 129
rect 1317 125 1318 129
rect 1312 123 1318 125
rect 1312 119 1313 123
rect 1317 119 1318 123
rect 1312 117 1318 119
rect 1312 113 1313 117
rect 1317 113 1318 117
rect 1312 111 1318 113
rect 1312 107 1313 111
rect 1317 107 1318 111
rect 1312 105 1318 107
rect 1312 101 1313 105
rect 1317 101 1318 105
rect 1312 99 1318 101
rect 1312 95 1313 99
rect 1317 95 1318 99
rect 1312 93 1318 95
rect 1312 89 1313 93
rect 1317 89 1318 93
rect 1312 87 1318 89
rect 1312 83 1313 87
rect 1317 83 1318 87
rect 1312 81 1318 83
rect 1312 77 1313 81
rect 1317 77 1318 81
rect 1312 75 1318 77
rect 1312 71 1313 75
rect 1317 71 1318 75
rect 1312 69 1318 71
rect 1312 65 1313 69
rect 1317 65 1318 69
rect 1312 63 1318 65
rect 1312 59 1313 63
rect 1317 59 1318 63
rect 1312 57 1318 59
rect 1312 53 1313 57
rect 1317 53 1318 57
rect 1312 51 1318 53
rect 1312 47 1313 51
rect 1317 47 1318 51
rect 1312 45 1318 47
rect 1312 41 1313 45
rect 1317 41 1318 45
rect 1312 39 1318 41
rect 1312 35 1313 39
rect 1317 35 1318 39
rect 1312 33 1318 35
rect 1312 29 1313 33
rect 1317 29 1318 33
rect 1312 27 1318 29
rect 1312 23 1313 27
rect 1317 23 1318 27
rect 1312 21 1318 23
rect 1312 17 1313 21
rect 1317 17 1318 21
rect 1312 15 1318 17
rect 1312 11 1313 15
rect 1317 11 1318 15
rect 1312 9 1318 11
rect 1312 5 1313 9
rect 1317 5 1318 9
rect 1312 2 1318 5
rect 1786 363 1792 364
rect 1786 359 1787 363
rect 1791 359 1792 363
rect 1786 357 1792 359
rect 1786 353 1787 357
rect 1791 353 1792 357
rect 1786 351 1792 353
rect 1786 347 1787 351
rect 1791 347 1792 351
rect 1786 345 1792 347
rect 1786 341 1787 345
rect 1791 341 1792 345
rect 1786 339 1792 341
rect 1786 335 1787 339
rect 1791 335 1792 339
rect 1786 333 1792 335
rect 1786 329 1787 333
rect 1791 329 1792 333
rect 1786 327 1792 329
rect 1786 323 1787 327
rect 1791 323 1792 327
rect 1786 321 1792 323
rect 1786 317 1787 321
rect 1791 317 1792 321
rect 1786 315 1792 317
rect 1786 311 1787 315
rect 1791 311 1792 315
rect 1786 309 1792 311
rect 1786 305 1787 309
rect 1791 305 1792 309
rect 1786 303 1792 305
rect 1786 299 1787 303
rect 1791 299 1792 303
rect 1786 297 1792 299
rect 1786 293 1787 297
rect 1791 293 1792 297
rect 1786 291 1792 293
rect 1786 287 1787 291
rect 1791 287 1792 291
rect 1786 285 1792 287
rect 1786 281 1787 285
rect 1791 281 1792 285
rect 1786 279 1792 281
rect 1786 275 1787 279
rect 1791 275 1792 279
rect 1786 273 1792 275
rect 1786 269 1787 273
rect 1791 269 1792 273
rect 1786 267 1792 269
rect 1786 263 1787 267
rect 1791 263 1792 267
rect 1786 261 1792 263
rect 1786 257 1787 261
rect 1791 257 1792 261
rect 1786 255 1792 257
rect 1786 251 1787 255
rect 1791 251 1792 255
rect 1786 249 1792 251
rect 1786 245 1787 249
rect 1791 245 1792 249
rect 1786 243 1792 245
rect 1786 239 1787 243
rect 1791 239 1792 243
rect 1786 237 1792 239
rect 1786 233 1787 237
rect 1791 233 1792 237
rect 1786 231 1792 233
rect 1786 227 1787 231
rect 1791 227 1792 231
rect 1786 225 1792 227
rect 1786 221 1787 225
rect 1791 221 1792 225
rect 1786 219 1792 221
rect 1786 215 1787 219
rect 1791 215 1792 219
rect 1786 213 1792 215
rect 1786 209 1787 213
rect 1791 209 1792 213
rect 1786 207 1792 209
rect 1786 203 1787 207
rect 1791 203 1792 207
rect 1786 201 1792 203
rect 1786 197 1787 201
rect 1791 197 1792 201
rect 1786 195 1792 197
rect 1786 191 1787 195
rect 1791 191 1792 195
rect 1786 189 1792 191
rect 1786 185 1787 189
rect 1791 185 1792 189
rect 1786 183 1792 185
rect 1786 179 1787 183
rect 1791 179 1792 183
rect 1786 177 1792 179
rect 1786 173 1787 177
rect 1791 173 1792 177
rect 1786 171 1792 173
rect 1786 167 1787 171
rect 1791 167 1792 171
rect 1786 165 1792 167
rect 1786 161 1787 165
rect 1791 161 1792 165
rect 1786 159 1792 161
rect 1786 155 1787 159
rect 1791 155 1792 159
rect 1786 153 1792 155
rect 1786 149 1787 153
rect 1791 149 1792 153
rect 1786 147 1792 149
rect 1786 143 1787 147
rect 1791 143 1792 147
rect 1786 141 1792 143
rect 1786 137 1787 141
rect 1791 137 1792 141
rect 1786 135 1792 137
rect 1786 131 1787 135
rect 1791 131 1792 135
rect 1786 129 1792 131
rect 1786 125 1787 129
rect 1791 125 1792 129
rect 1786 123 1792 125
rect 1786 119 1787 123
rect 1791 119 1792 123
rect 1786 117 1792 119
rect 1786 113 1787 117
rect 1791 113 1792 117
rect 1786 111 1792 113
rect 1786 107 1787 111
rect 1791 107 1792 111
rect 1786 105 1792 107
rect 1786 101 1787 105
rect 1791 101 1792 105
rect 1786 99 1792 101
rect 1786 95 1787 99
rect 1791 95 1792 99
rect 1786 93 1792 95
rect 1786 89 1787 93
rect 1791 89 1792 93
rect 1786 87 1792 89
rect 1786 83 1787 87
rect 1791 83 1792 87
rect 1786 81 1792 83
rect 1786 77 1787 81
rect 1791 77 1792 81
rect 1786 75 1792 77
rect 1786 71 1787 75
rect 1791 71 1792 75
rect 1786 69 1792 71
rect 1786 65 1787 69
rect 1791 65 1792 69
rect 1786 63 1792 65
rect 1786 59 1787 63
rect 1791 59 1792 63
rect 1786 57 1792 59
rect 1786 53 1787 57
rect 1791 53 1792 57
rect 1786 51 1792 53
rect 1786 47 1787 51
rect 1791 47 1792 51
rect 1786 45 1792 47
rect 1786 41 1787 45
rect 1791 41 1792 45
rect 1786 39 1792 41
rect 1786 35 1787 39
rect 1791 35 1792 39
rect 1786 33 1792 35
rect 1786 29 1787 33
rect 1791 29 1792 33
rect 1786 27 1792 29
rect 1786 23 1787 27
rect 1791 23 1792 27
rect 1786 21 1792 23
rect 1786 17 1787 21
rect 1791 17 1792 21
rect 1786 15 1792 17
rect 1786 11 1787 15
rect 1791 11 1792 15
rect 1786 9 1792 11
rect 1786 5 1787 9
rect 1791 5 1792 9
rect 1786 2 1792 5
rect 2260 363 2266 364
rect 2260 359 2261 363
rect 2265 359 2266 363
rect 2260 357 2266 359
rect 2260 353 2261 357
rect 2265 353 2266 357
rect 2260 351 2266 353
rect 2260 347 2261 351
rect 2265 347 2266 351
rect 2260 345 2266 347
rect 2260 341 2261 345
rect 2265 341 2266 345
rect 2260 339 2266 341
rect 2260 335 2261 339
rect 2265 335 2266 339
rect 2260 333 2266 335
rect 2260 329 2261 333
rect 2265 329 2266 333
rect 2260 327 2266 329
rect 2260 323 2261 327
rect 2265 323 2266 327
rect 2260 321 2266 323
rect 2260 317 2261 321
rect 2265 317 2266 321
rect 2260 315 2266 317
rect 2260 311 2261 315
rect 2265 311 2266 315
rect 2260 309 2266 311
rect 2260 305 2261 309
rect 2265 305 2266 309
rect 2260 303 2266 305
rect 2260 299 2261 303
rect 2265 299 2266 303
rect 2260 297 2266 299
rect 2260 293 2261 297
rect 2265 293 2266 297
rect 2260 291 2266 293
rect 2260 287 2261 291
rect 2265 287 2266 291
rect 2260 285 2266 287
rect 2260 281 2261 285
rect 2265 281 2266 285
rect 2260 279 2266 281
rect 2260 275 2261 279
rect 2265 275 2266 279
rect 2260 273 2266 275
rect 2260 269 2261 273
rect 2265 269 2266 273
rect 2260 267 2266 269
rect 2260 263 2261 267
rect 2265 263 2266 267
rect 2260 261 2266 263
rect 2260 257 2261 261
rect 2265 257 2266 261
rect 2260 255 2266 257
rect 2260 251 2261 255
rect 2265 251 2266 255
rect 2260 249 2266 251
rect 2260 245 2261 249
rect 2265 245 2266 249
rect 2260 243 2266 245
rect 2260 239 2261 243
rect 2265 239 2266 243
rect 2260 237 2266 239
rect 2260 233 2261 237
rect 2265 233 2266 237
rect 2260 231 2266 233
rect 2260 227 2261 231
rect 2265 227 2266 231
rect 2260 225 2266 227
rect 2260 221 2261 225
rect 2265 221 2266 225
rect 2260 219 2266 221
rect 2260 215 2261 219
rect 2265 215 2266 219
rect 2260 213 2266 215
rect 2260 209 2261 213
rect 2265 209 2266 213
rect 2260 207 2266 209
rect 2260 203 2261 207
rect 2265 203 2266 207
rect 2260 201 2266 203
rect 2260 197 2261 201
rect 2265 197 2266 201
rect 2260 195 2266 197
rect 2260 191 2261 195
rect 2265 191 2266 195
rect 2260 189 2266 191
rect 2260 185 2261 189
rect 2265 185 2266 189
rect 2260 183 2266 185
rect 2260 179 2261 183
rect 2265 179 2266 183
rect 2260 177 2266 179
rect 2260 173 2261 177
rect 2265 173 2266 177
rect 2260 171 2266 173
rect 2260 167 2261 171
rect 2265 167 2266 171
rect 2260 165 2266 167
rect 2260 161 2261 165
rect 2265 161 2266 165
rect 2260 159 2266 161
rect 2260 155 2261 159
rect 2265 155 2266 159
rect 2260 153 2266 155
rect 2260 149 2261 153
rect 2265 149 2266 153
rect 2260 147 2266 149
rect 2260 143 2261 147
rect 2265 143 2266 147
rect 2260 141 2266 143
rect 2260 137 2261 141
rect 2265 137 2266 141
rect 2260 135 2266 137
rect 2260 131 2261 135
rect 2265 131 2266 135
rect 2260 129 2266 131
rect 2260 125 2261 129
rect 2265 125 2266 129
rect 2260 123 2266 125
rect 2260 119 2261 123
rect 2265 119 2266 123
rect 2260 117 2266 119
rect 2260 113 2261 117
rect 2265 113 2266 117
rect 2260 111 2266 113
rect 2260 107 2261 111
rect 2265 107 2266 111
rect 2260 105 2266 107
rect 2260 101 2261 105
rect 2265 101 2266 105
rect 2260 99 2266 101
rect 2260 95 2261 99
rect 2265 95 2266 99
rect 2260 93 2266 95
rect 2260 89 2261 93
rect 2265 89 2266 93
rect 2260 87 2266 89
rect 2260 83 2261 87
rect 2265 83 2266 87
rect 2260 81 2266 83
rect 2260 77 2261 81
rect 2265 77 2266 81
rect 2260 75 2266 77
rect 2260 71 2261 75
rect 2265 71 2266 75
rect 2260 69 2266 71
rect 2260 65 2261 69
rect 2265 65 2266 69
rect 2260 63 2266 65
rect 2260 59 2261 63
rect 2265 59 2266 63
rect 2260 57 2266 59
rect 2260 53 2261 57
rect 2265 53 2266 57
rect 2260 51 2266 53
rect 2260 47 2261 51
rect 2265 47 2266 51
rect 2260 45 2266 47
rect 2260 41 2261 45
rect 2265 41 2266 45
rect 2260 39 2266 41
rect 2260 35 2261 39
rect 2265 35 2266 39
rect 2260 33 2266 35
rect 2260 29 2261 33
rect 2265 29 2266 33
rect 2260 27 2266 29
rect 2260 23 2261 27
rect 2265 23 2266 27
rect 2260 21 2266 23
rect 2260 17 2261 21
rect 2265 17 2266 21
rect 2260 15 2266 17
rect 2260 11 2261 15
rect 2265 11 2266 15
rect 2260 9 2266 11
rect 2260 5 2261 9
rect 2265 5 2266 9
rect 2260 2 2266 5
rect 2734 363 2740 364
rect 2734 359 2735 363
rect 2739 359 2740 363
rect 2734 357 2740 359
rect 2734 353 2735 357
rect 2739 353 2740 357
rect 2734 351 2740 353
rect 2734 347 2735 351
rect 2739 347 2740 351
rect 2734 345 2740 347
rect 2734 341 2735 345
rect 2739 341 2740 345
rect 2734 339 2740 341
rect 2734 335 2735 339
rect 2739 335 2740 339
rect 2734 333 2740 335
rect 2734 329 2735 333
rect 2739 329 2740 333
rect 2734 327 2740 329
rect 2734 323 2735 327
rect 2739 323 2740 327
rect 2734 321 2740 323
rect 2734 317 2735 321
rect 2739 317 2740 321
rect 2734 315 2740 317
rect 2734 311 2735 315
rect 2739 311 2740 315
rect 2734 309 2740 311
rect 2734 305 2735 309
rect 2739 305 2740 309
rect 2734 303 2740 305
rect 2734 299 2735 303
rect 2739 299 2740 303
rect 2734 297 2740 299
rect 2734 293 2735 297
rect 2739 293 2740 297
rect 2734 291 2740 293
rect 2734 287 2735 291
rect 2739 287 2740 291
rect 2734 285 2740 287
rect 2734 281 2735 285
rect 2739 281 2740 285
rect 2734 279 2740 281
rect 2734 275 2735 279
rect 2739 275 2740 279
rect 2734 273 2740 275
rect 2734 269 2735 273
rect 2739 269 2740 273
rect 2734 267 2740 269
rect 2734 263 2735 267
rect 2739 263 2740 267
rect 2734 261 2740 263
rect 2734 257 2735 261
rect 2739 257 2740 261
rect 2734 255 2740 257
rect 2734 251 2735 255
rect 2739 251 2740 255
rect 2734 249 2740 251
rect 2734 245 2735 249
rect 2739 245 2740 249
rect 2734 243 2740 245
rect 2734 239 2735 243
rect 2739 239 2740 243
rect 2734 237 2740 239
rect 2734 233 2735 237
rect 2739 233 2740 237
rect 2734 231 2740 233
rect 2734 227 2735 231
rect 2739 227 2740 231
rect 2734 225 2740 227
rect 2734 221 2735 225
rect 2739 221 2740 225
rect 2734 219 2740 221
rect 2734 215 2735 219
rect 2739 215 2740 219
rect 2734 213 2740 215
rect 2734 209 2735 213
rect 2739 209 2740 213
rect 2734 207 2740 209
rect 2734 203 2735 207
rect 2739 203 2740 207
rect 2734 201 2740 203
rect 2734 197 2735 201
rect 2739 197 2740 201
rect 2734 195 2740 197
rect 2734 191 2735 195
rect 2739 191 2740 195
rect 2734 189 2740 191
rect 2734 185 2735 189
rect 2739 185 2740 189
rect 2734 183 2740 185
rect 2734 179 2735 183
rect 2739 179 2740 183
rect 2734 177 2740 179
rect 2734 173 2735 177
rect 2739 173 2740 177
rect 2734 171 2740 173
rect 2734 167 2735 171
rect 2739 167 2740 171
rect 2734 165 2740 167
rect 2734 161 2735 165
rect 2739 161 2740 165
rect 2734 159 2740 161
rect 2734 155 2735 159
rect 2739 155 2740 159
rect 2734 153 2740 155
rect 2734 149 2735 153
rect 2739 149 2740 153
rect 2734 147 2740 149
rect 2734 143 2735 147
rect 2739 143 2740 147
rect 2734 141 2740 143
rect 2734 137 2735 141
rect 2739 137 2740 141
rect 2734 135 2740 137
rect 2734 131 2735 135
rect 2739 131 2740 135
rect 2734 129 2740 131
rect 2734 125 2735 129
rect 2739 125 2740 129
rect 2734 123 2740 125
rect 2734 119 2735 123
rect 2739 119 2740 123
rect 2734 117 2740 119
rect 2734 113 2735 117
rect 2739 113 2740 117
rect 2734 111 2740 113
rect 2734 107 2735 111
rect 2739 107 2740 111
rect 2734 105 2740 107
rect 2734 101 2735 105
rect 2739 101 2740 105
rect 2734 99 2740 101
rect 2734 95 2735 99
rect 2739 95 2740 99
rect 2734 93 2740 95
rect 2734 89 2735 93
rect 2739 89 2740 93
rect 2734 87 2740 89
rect 2734 83 2735 87
rect 2739 83 2740 87
rect 2734 81 2740 83
rect 2734 77 2735 81
rect 2739 77 2740 81
rect 2734 75 2740 77
rect 2734 71 2735 75
rect 2739 71 2740 75
rect 2734 69 2740 71
rect 2734 65 2735 69
rect 2739 65 2740 69
rect 2734 63 2740 65
rect 2734 59 2735 63
rect 2739 59 2740 63
rect 2734 57 2740 59
rect 2734 53 2735 57
rect 2739 53 2740 57
rect 2734 51 2740 53
rect 2734 47 2735 51
rect 2739 47 2740 51
rect 2734 45 2740 47
rect 2734 41 2735 45
rect 2739 41 2740 45
rect 2734 39 2740 41
rect 2734 35 2735 39
rect 2739 35 2740 39
rect 2734 33 2740 35
rect 2734 29 2735 33
rect 2739 29 2740 33
rect 2734 27 2740 29
rect 2734 23 2735 27
rect 2739 23 2740 27
rect 2734 21 2740 23
rect 2734 17 2735 21
rect 2739 17 2740 21
rect 2734 15 2740 17
rect 2734 11 2735 15
rect 2739 11 2740 15
rect 2734 9 2740 11
rect 2734 5 2735 9
rect 2739 5 2740 9
rect 2734 2 2740 5
rect 3208 363 3214 364
rect 3208 359 3209 363
rect 3213 359 3214 363
rect 3208 357 3214 359
rect 3208 353 3209 357
rect 3213 353 3214 357
rect 3208 351 3214 353
rect 3208 347 3209 351
rect 3213 347 3214 351
rect 3208 345 3214 347
rect 3208 341 3209 345
rect 3213 341 3214 345
rect 3208 339 3214 341
rect 3208 335 3209 339
rect 3213 335 3214 339
rect 3208 333 3214 335
rect 3208 329 3209 333
rect 3213 329 3214 333
rect 3208 327 3214 329
rect 3208 323 3209 327
rect 3213 323 3214 327
rect 3208 321 3214 323
rect 3208 317 3209 321
rect 3213 317 3214 321
rect 3208 315 3214 317
rect 3208 311 3209 315
rect 3213 311 3214 315
rect 3208 309 3214 311
rect 3208 305 3209 309
rect 3213 305 3214 309
rect 3208 303 3214 305
rect 3208 299 3209 303
rect 3213 299 3214 303
rect 3208 297 3214 299
rect 3208 293 3209 297
rect 3213 293 3214 297
rect 3208 291 3214 293
rect 3208 287 3209 291
rect 3213 287 3214 291
rect 3208 285 3214 287
rect 3208 281 3209 285
rect 3213 281 3214 285
rect 3208 279 3214 281
rect 3208 275 3209 279
rect 3213 275 3214 279
rect 3208 273 3214 275
rect 3208 269 3209 273
rect 3213 269 3214 273
rect 3208 267 3214 269
rect 3208 263 3209 267
rect 3213 263 3214 267
rect 3208 261 3214 263
rect 3208 257 3209 261
rect 3213 257 3214 261
rect 3208 255 3214 257
rect 3208 251 3209 255
rect 3213 251 3214 255
rect 3208 249 3214 251
rect 3208 245 3209 249
rect 3213 245 3214 249
rect 3208 243 3214 245
rect 3208 239 3209 243
rect 3213 239 3214 243
rect 3208 237 3214 239
rect 3208 233 3209 237
rect 3213 233 3214 237
rect 3208 231 3214 233
rect 3208 227 3209 231
rect 3213 227 3214 231
rect 3208 225 3214 227
rect 3208 221 3209 225
rect 3213 221 3214 225
rect 3208 219 3214 221
rect 3208 215 3209 219
rect 3213 215 3214 219
rect 3208 213 3214 215
rect 3208 209 3209 213
rect 3213 209 3214 213
rect 3208 207 3214 209
rect 3208 203 3209 207
rect 3213 203 3214 207
rect 3208 201 3214 203
rect 3208 197 3209 201
rect 3213 197 3214 201
rect 3208 195 3214 197
rect 3208 191 3209 195
rect 3213 191 3214 195
rect 3208 189 3214 191
rect 3208 185 3209 189
rect 3213 185 3214 189
rect 3208 183 3214 185
rect 3208 179 3209 183
rect 3213 179 3214 183
rect 3208 177 3214 179
rect 3208 173 3209 177
rect 3213 173 3214 177
rect 3208 171 3214 173
rect 3208 167 3209 171
rect 3213 167 3214 171
rect 3208 165 3214 167
rect 3208 161 3209 165
rect 3213 161 3214 165
rect 3208 159 3214 161
rect 3208 155 3209 159
rect 3213 155 3214 159
rect 3208 153 3214 155
rect 3208 149 3209 153
rect 3213 149 3214 153
rect 3208 147 3214 149
rect 3208 143 3209 147
rect 3213 143 3214 147
rect 3208 141 3214 143
rect 3208 137 3209 141
rect 3213 137 3214 141
rect 3208 135 3214 137
rect 3208 131 3209 135
rect 3213 131 3214 135
rect 3208 129 3214 131
rect 3208 125 3209 129
rect 3213 125 3214 129
rect 3208 123 3214 125
rect 3208 119 3209 123
rect 3213 119 3214 123
rect 3208 117 3214 119
rect 3208 113 3209 117
rect 3213 113 3214 117
rect 3208 111 3214 113
rect 3208 107 3209 111
rect 3213 107 3214 111
rect 3208 105 3214 107
rect 3208 101 3209 105
rect 3213 101 3214 105
rect 3208 99 3214 101
rect 3208 95 3209 99
rect 3213 95 3214 99
rect 3208 93 3214 95
rect 3208 89 3209 93
rect 3213 89 3214 93
rect 3208 87 3214 89
rect 3208 83 3209 87
rect 3213 83 3214 87
rect 3208 81 3214 83
rect 3208 77 3209 81
rect 3213 77 3214 81
rect 3208 75 3214 77
rect 3208 71 3209 75
rect 3213 71 3214 75
rect 3208 69 3214 71
rect 3208 65 3209 69
rect 3213 65 3214 69
rect 3208 63 3214 65
rect 3208 59 3209 63
rect 3213 59 3214 63
rect 3208 57 3214 59
rect 3208 53 3209 57
rect 3213 53 3214 57
rect 3208 51 3214 53
rect 3208 47 3209 51
rect 3213 47 3214 51
rect 3208 45 3214 47
rect 3208 41 3209 45
rect 3213 41 3214 45
rect 3208 39 3214 41
rect 3208 35 3209 39
rect 3213 35 3214 39
rect 3208 33 3214 35
rect 3208 29 3209 33
rect 3213 29 3214 33
rect 3208 27 3214 29
rect 3208 23 3209 27
rect 3213 23 3214 27
rect 3208 21 3214 23
rect 3208 17 3209 21
rect 3213 17 3214 21
rect 3208 15 3214 17
rect 3208 11 3209 15
rect 3213 11 3214 15
rect 3208 9 3214 11
rect 3208 5 3209 9
rect 3213 5 3214 9
rect 3208 2 3214 5
rect 3682 363 3688 364
rect 3682 359 3683 363
rect 3687 359 3688 363
rect 3682 357 3688 359
rect 3682 353 3683 357
rect 3687 353 3688 357
rect 3682 351 3688 353
rect 3682 347 3683 351
rect 3687 347 3688 351
rect 3682 345 3688 347
rect 3682 341 3683 345
rect 3687 341 3688 345
rect 3682 339 3688 341
rect 3682 335 3683 339
rect 3687 335 3688 339
rect 3682 333 3688 335
rect 3682 329 3683 333
rect 3687 329 3688 333
rect 3682 327 3688 329
rect 3682 323 3683 327
rect 3687 323 3688 327
rect 3682 321 3688 323
rect 3682 317 3683 321
rect 3687 317 3688 321
rect 3682 315 3688 317
rect 3682 311 3683 315
rect 3687 311 3688 315
rect 3682 309 3688 311
rect 3682 305 3683 309
rect 3687 305 3688 309
rect 3682 303 3688 305
rect 3682 299 3683 303
rect 3687 299 3688 303
rect 3682 297 3688 299
rect 3682 293 3683 297
rect 3687 293 3688 297
rect 3682 291 3688 293
rect 3682 287 3683 291
rect 3687 287 3688 291
rect 3682 285 3688 287
rect 3682 281 3683 285
rect 3687 281 3688 285
rect 3682 279 3688 281
rect 3682 275 3683 279
rect 3687 275 3688 279
rect 3682 273 3688 275
rect 3682 269 3683 273
rect 3687 269 3688 273
rect 3682 267 3688 269
rect 3682 263 3683 267
rect 3687 263 3688 267
rect 3682 261 3688 263
rect 3682 257 3683 261
rect 3687 257 3688 261
rect 3682 255 3688 257
rect 3682 251 3683 255
rect 3687 251 3688 255
rect 3682 249 3688 251
rect 3682 245 3683 249
rect 3687 245 3688 249
rect 3682 243 3688 245
rect 3682 239 3683 243
rect 3687 239 3688 243
rect 3682 237 3688 239
rect 3682 233 3683 237
rect 3687 233 3688 237
rect 3682 231 3688 233
rect 3682 227 3683 231
rect 3687 227 3688 231
rect 3682 225 3688 227
rect 3682 221 3683 225
rect 3687 221 3688 225
rect 3682 219 3688 221
rect 3682 215 3683 219
rect 3687 215 3688 219
rect 3682 213 3688 215
rect 3682 209 3683 213
rect 3687 209 3688 213
rect 3682 207 3688 209
rect 3682 203 3683 207
rect 3687 203 3688 207
rect 3682 201 3688 203
rect 3682 197 3683 201
rect 3687 197 3688 201
rect 3682 195 3688 197
rect 3682 191 3683 195
rect 3687 191 3688 195
rect 3682 189 3688 191
rect 3682 185 3683 189
rect 3687 185 3688 189
rect 3682 183 3688 185
rect 3682 179 3683 183
rect 3687 179 3688 183
rect 3682 177 3688 179
rect 3682 173 3683 177
rect 3687 173 3688 177
rect 3682 171 3688 173
rect 3682 167 3683 171
rect 3687 167 3688 171
rect 3682 165 3688 167
rect 3682 161 3683 165
rect 3687 161 3688 165
rect 3682 159 3688 161
rect 3682 155 3683 159
rect 3687 155 3688 159
rect 3682 153 3688 155
rect 3682 149 3683 153
rect 3687 149 3688 153
rect 3682 147 3688 149
rect 3682 143 3683 147
rect 3687 143 3688 147
rect 3682 141 3688 143
rect 3682 137 3683 141
rect 3687 137 3688 141
rect 3682 135 3688 137
rect 3682 131 3683 135
rect 3687 131 3688 135
rect 3682 129 3688 131
rect 3682 125 3683 129
rect 3687 125 3688 129
rect 3682 123 3688 125
rect 3682 119 3683 123
rect 3687 119 3688 123
rect 3682 117 3688 119
rect 3682 113 3683 117
rect 3687 113 3688 117
rect 3682 111 3688 113
rect 3682 107 3683 111
rect 3687 107 3688 111
rect 3682 105 3688 107
rect 3682 101 3683 105
rect 3687 101 3688 105
rect 3682 99 3688 101
rect 3682 95 3683 99
rect 3687 95 3688 99
rect 3682 93 3688 95
rect 3682 89 3683 93
rect 3687 89 3688 93
rect 3682 87 3688 89
rect 3682 83 3683 87
rect 3687 83 3688 87
rect 3682 81 3688 83
rect 3682 77 3683 81
rect 3687 77 3688 81
rect 3682 75 3688 77
rect 3682 71 3683 75
rect 3687 71 3688 75
rect 3682 69 3688 71
rect 3682 65 3683 69
rect 3687 65 3688 69
rect 3682 63 3688 65
rect 3682 59 3683 63
rect 3687 59 3688 63
rect 3682 57 3688 59
rect 3682 53 3683 57
rect 3687 53 3688 57
rect 3682 51 3688 53
rect 3682 47 3683 51
rect 3687 47 3688 51
rect 3682 45 3688 47
rect 3682 41 3683 45
rect 3687 41 3688 45
rect 3682 39 3688 41
rect 3682 35 3683 39
rect 3687 35 3688 39
rect 3682 33 3688 35
rect 3682 29 3683 33
rect 3687 29 3688 33
rect 3682 27 3688 29
rect 3682 23 3683 27
rect 3687 23 3688 27
rect 3682 21 3688 23
rect 3682 17 3683 21
rect 3687 17 3688 21
rect 3682 15 3688 17
rect 3682 11 3683 15
rect 3687 11 3688 15
rect 3682 9 3688 11
rect 3682 5 3683 9
rect 3687 5 3688 9
rect 3682 2 3688 5
rect 4156 363 4162 364
rect 4156 359 4157 363
rect 4161 359 4162 363
rect 4156 357 4162 359
rect 4156 353 4157 357
rect 4161 353 4162 357
rect 4156 351 4162 353
rect 4156 347 4157 351
rect 4161 347 4162 351
rect 4156 345 4162 347
rect 4156 341 4157 345
rect 4161 341 4162 345
rect 4156 339 4162 341
rect 4156 335 4157 339
rect 4161 335 4162 339
rect 4156 333 4162 335
rect 4156 329 4157 333
rect 4161 329 4162 333
rect 4156 327 4162 329
rect 4156 323 4157 327
rect 4161 323 4162 327
rect 4156 321 4162 323
rect 4156 317 4157 321
rect 4161 317 4162 321
rect 4156 315 4162 317
rect 4156 311 4157 315
rect 4161 311 4162 315
rect 4156 309 4162 311
rect 4156 305 4157 309
rect 4161 305 4162 309
rect 4156 303 4162 305
rect 4156 299 4157 303
rect 4161 299 4162 303
rect 4156 297 4162 299
rect 4156 293 4157 297
rect 4161 293 4162 297
rect 4156 291 4162 293
rect 4156 287 4157 291
rect 4161 287 4162 291
rect 4156 285 4162 287
rect 4156 281 4157 285
rect 4161 281 4162 285
rect 4156 279 4162 281
rect 4156 275 4157 279
rect 4161 275 4162 279
rect 4156 273 4162 275
rect 4156 269 4157 273
rect 4161 269 4162 273
rect 4156 267 4162 269
rect 4156 263 4157 267
rect 4161 263 4162 267
rect 4156 261 4162 263
rect 4156 257 4157 261
rect 4161 257 4162 261
rect 4156 255 4162 257
rect 4156 251 4157 255
rect 4161 251 4162 255
rect 4156 249 4162 251
rect 4156 245 4157 249
rect 4161 245 4162 249
rect 4156 243 4162 245
rect 4156 239 4157 243
rect 4161 239 4162 243
rect 4156 237 4162 239
rect 4156 233 4157 237
rect 4161 233 4162 237
rect 4156 231 4162 233
rect 4156 227 4157 231
rect 4161 227 4162 231
rect 4156 225 4162 227
rect 4156 221 4157 225
rect 4161 221 4162 225
rect 4156 219 4162 221
rect 4156 215 4157 219
rect 4161 215 4162 219
rect 4156 213 4162 215
rect 4156 209 4157 213
rect 4161 209 4162 213
rect 4156 207 4162 209
rect 4156 203 4157 207
rect 4161 203 4162 207
rect 4156 201 4162 203
rect 4156 197 4157 201
rect 4161 197 4162 201
rect 4156 195 4162 197
rect 4156 191 4157 195
rect 4161 191 4162 195
rect 4156 189 4162 191
rect 4156 185 4157 189
rect 4161 185 4162 189
rect 4156 183 4162 185
rect 4156 179 4157 183
rect 4161 179 4162 183
rect 4156 177 4162 179
rect 4156 173 4157 177
rect 4161 173 4162 177
rect 4156 171 4162 173
rect 4156 167 4157 171
rect 4161 167 4162 171
rect 4156 165 4162 167
rect 4156 161 4157 165
rect 4161 161 4162 165
rect 4156 159 4162 161
rect 4156 155 4157 159
rect 4161 155 4162 159
rect 4156 153 4162 155
rect 4156 149 4157 153
rect 4161 149 4162 153
rect 4156 147 4162 149
rect 4156 143 4157 147
rect 4161 143 4162 147
rect 4156 141 4162 143
rect 4156 137 4157 141
rect 4161 137 4162 141
rect 4156 135 4162 137
rect 4156 131 4157 135
rect 4161 131 4162 135
rect 4156 129 4162 131
rect 4156 125 4157 129
rect 4161 125 4162 129
rect 4156 123 4162 125
rect 4156 119 4157 123
rect 4161 119 4162 123
rect 4156 117 4162 119
rect 4156 113 4157 117
rect 4161 113 4162 117
rect 4156 111 4162 113
rect 4156 107 4157 111
rect 4161 107 4162 111
rect 4156 105 4162 107
rect 4156 101 4157 105
rect 4161 101 4162 105
rect 4156 99 4162 101
rect 4156 95 4157 99
rect 4161 95 4162 99
rect 4156 93 4162 95
rect 4156 89 4157 93
rect 4161 89 4162 93
rect 4156 87 4162 89
rect 4156 83 4157 87
rect 4161 83 4162 87
rect 4156 81 4162 83
rect 4156 77 4157 81
rect 4161 77 4162 81
rect 4156 75 4162 77
rect 4156 71 4157 75
rect 4161 71 4162 75
rect 4156 69 4162 71
rect 4156 65 4157 69
rect 4161 65 4162 69
rect 4156 63 4162 65
rect 4156 59 4157 63
rect 4161 59 4162 63
rect 4156 57 4162 59
rect 4156 53 4157 57
rect 4161 53 4162 57
rect 4156 51 4162 53
rect 4156 47 4157 51
rect 4161 47 4162 51
rect 4156 45 4162 47
rect 4156 41 4157 45
rect 4161 41 4162 45
rect 4156 39 4162 41
rect 4156 35 4157 39
rect 4161 35 4162 39
rect 4156 33 4162 35
rect 4156 29 4157 33
rect 4161 29 4162 33
rect 4156 27 4162 29
rect 4156 23 4157 27
rect 4161 23 4162 27
rect 4156 21 4162 23
rect 4156 17 4157 21
rect 4161 17 4162 21
rect 4156 15 4162 17
rect 4156 11 4157 15
rect 4161 11 4162 15
rect 4156 9 4162 11
rect 4156 5 4157 9
rect 4161 5 4162 9
rect 4156 2 4162 5
rect 4630 363 4636 364
rect 4630 359 4631 363
rect 4635 359 4636 363
rect 4630 357 4636 359
rect 4630 353 4631 357
rect 4635 353 4636 357
rect 4630 351 4636 353
rect 4630 347 4631 351
rect 4635 347 4636 351
rect 4630 345 4636 347
rect 4630 341 4631 345
rect 4635 341 4636 345
rect 4630 339 4636 341
rect 4630 335 4631 339
rect 4635 335 4636 339
rect 4630 333 4636 335
rect 4630 329 4631 333
rect 4635 329 4636 333
rect 4630 327 4636 329
rect 4630 323 4631 327
rect 4635 323 4636 327
rect 4630 321 4636 323
rect 4630 317 4631 321
rect 4635 317 4636 321
rect 4630 315 4636 317
rect 4630 311 4631 315
rect 4635 311 4636 315
rect 4630 309 4636 311
rect 4630 305 4631 309
rect 4635 305 4636 309
rect 4630 303 4636 305
rect 4630 299 4631 303
rect 4635 299 4636 303
rect 4630 297 4636 299
rect 4630 293 4631 297
rect 4635 293 4636 297
rect 4630 291 4636 293
rect 4630 287 4631 291
rect 4635 287 4636 291
rect 4630 285 4636 287
rect 4630 281 4631 285
rect 4635 281 4636 285
rect 4630 279 4636 281
rect 4630 275 4631 279
rect 4635 275 4636 279
rect 4630 273 4636 275
rect 4630 269 4631 273
rect 4635 269 4636 273
rect 4630 267 4636 269
rect 4630 263 4631 267
rect 4635 263 4636 267
rect 4630 261 4636 263
rect 4630 257 4631 261
rect 4635 257 4636 261
rect 4630 255 4636 257
rect 4630 251 4631 255
rect 4635 251 4636 255
rect 4630 249 4636 251
rect 4630 245 4631 249
rect 4635 245 4636 249
rect 4630 243 4636 245
rect 4630 239 4631 243
rect 4635 239 4636 243
rect 4630 237 4636 239
rect 4630 233 4631 237
rect 4635 233 4636 237
rect 4630 231 4636 233
rect 4630 227 4631 231
rect 4635 227 4636 231
rect 4630 225 4636 227
rect 4630 221 4631 225
rect 4635 221 4636 225
rect 4630 219 4636 221
rect 4630 215 4631 219
rect 4635 215 4636 219
rect 4630 213 4636 215
rect 4630 209 4631 213
rect 4635 209 4636 213
rect 4630 207 4636 209
rect 4630 203 4631 207
rect 4635 203 4636 207
rect 4630 201 4636 203
rect 4630 197 4631 201
rect 4635 197 4636 201
rect 4630 195 4636 197
rect 4630 191 4631 195
rect 4635 191 4636 195
rect 4630 189 4636 191
rect 4630 185 4631 189
rect 4635 185 4636 189
rect 4630 183 4636 185
rect 4630 179 4631 183
rect 4635 179 4636 183
rect 4630 177 4636 179
rect 4630 173 4631 177
rect 4635 173 4636 177
rect 4630 171 4636 173
rect 4630 167 4631 171
rect 4635 167 4636 171
rect 4630 165 4636 167
rect 4630 161 4631 165
rect 4635 161 4636 165
rect 4630 159 4636 161
rect 4630 155 4631 159
rect 4635 155 4636 159
rect 4630 153 4636 155
rect 4630 149 4631 153
rect 4635 149 4636 153
rect 4630 147 4636 149
rect 4630 143 4631 147
rect 4635 143 4636 147
rect 4630 141 4636 143
rect 4630 137 4631 141
rect 4635 137 4636 141
rect 4630 135 4636 137
rect 4630 131 4631 135
rect 4635 131 4636 135
rect 4630 129 4636 131
rect 4630 125 4631 129
rect 4635 125 4636 129
rect 4630 123 4636 125
rect 4630 119 4631 123
rect 4635 119 4636 123
rect 4630 117 4636 119
rect 4630 113 4631 117
rect 4635 113 4636 117
rect 4630 111 4636 113
rect 4630 107 4631 111
rect 4635 107 4636 111
rect 4630 105 4636 107
rect 4630 101 4631 105
rect 4635 101 4636 105
rect 4630 99 4636 101
rect 4630 95 4631 99
rect 4635 95 4636 99
rect 4630 93 4636 95
rect 4630 89 4631 93
rect 4635 89 4636 93
rect 4630 87 4636 89
rect 4630 83 4631 87
rect 4635 83 4636 87
rect 4630 81 4636 83
rect 4630 77 4631 81
rect 4635 77 4636 81
rect 4630 75 4636 77
rect 4630 71 4631 75
rect 4635 71 4636 75
rect 4630 69 4636 71
rect 4630 65 4631 69
rect 4635 65 4636 69
rect 4630 63 4636 65
rect 4630 59 4631 63
rect 4635 59 4636 63
rect 4630 57 4636 59
rect 4630 53 4631 57
rect 4635 53 4636 57
rect 4630 51 4636 53
rect 4630 47 4631 51
rect 4635 47 4636 51
rect 4630 45 4636 47
rect 4630 41 4631 45
rect 4635 41 4636 45
rect 4630 39 4636 41
rect 4630 35 4631 39
rect 4635 35 4636 39
rect 4630 33 4636 35
rect 4630 29 4631 33
rect 4635 29 4636 33
rect 4630 27 4636 29
rect 4630 23 4631 27
rect 4635 23 4636 27
rect 4630 21 4636 23
rect 4630 17 4631 21
rect 4635 17 4636 21
rect 4630 15 4636 17
rect 4630 11 4631 15
rect 4635 11 4636 15
rect 4630 9 4636 11
rect 4630 5 4631 9
rect 4635 5 4636 9
rect 4630 2 4636 5
<< psubstratepcontact >>
rect 5 365 9 369
rect 11 365 15 369
rect 17 365 21 369
rect 23 365 27 369
rect 29 365 33 369
rect 35 365 39 369
rect 41 365 45 369
rect 47 365 51 369
rect 53 365 57 369
rect 59 365 63 369
rect 65 365 69 369
rect 71 365 75 369
rect 77 365 81 369
rect 83 365 87 369
rect 89 365 93 369
rect 95 365 99 369
rect 101 365 105 369
rect 107 365 111 369
rect 113 365 117 369
rect 119 365 123 369
rect 125 365 129 369
rect 131 365 135 369
rect 137 365 141 369
rect 143 365 147 369
rect 149 365 153 369
rect 155 365 159 369
rect 161 365 165 369
rect 167 365 171 369
rect 173 365 177 369
rect 179 365 183 369
rect 185 365 189 369
rect 191 365 195 369
rect 197 365 201 369
rect 203 365 207 369
rect 209 365 213 369
rect 215 365 219 369
rect 221 365 225 369
rect 227 365 231 369
rect 233 365 237 369
rect 239 365 243 369
rect 245 365 249 369
rect 251 365 255 369
rect 257 365 261 369
rect 263 365 267 369
rect 269 365 273 369
rect 275 365 279 369
rect 281 365 285 369
rect 287 365 291 369
rect 293 365 297 369
rect 299 365 303 369
rect 305 365 309 369
rect 311 365 315 369
rect 317 365 321 369
rect 323 365 327 369
rect 329 365 333 369
rect 335 365 339 369
rect 341 365 345 369
rect 347 365 351 369
rect 353 365 357 369
rect 359 365 363 369
rect 365 365 369 369
rect 371 365 375 369
rect 377 365 381 369
rect 383 365 387 369
rect 389 365 393 369
rect 395 365 399 369
rect 401 365 405 369
rect 407 365 411 369
rect 413 365 417 369
rect 419 365 423 369
rect 425 365 429 369
rect 431 365 435 369
rect 437 365 441 369
rect 443 365 447 369
rect 449 365 453 369
rect 455 365 459 369
rect 461 365 465 369
rect 467 365 471 369
rect 473 365 477 369
rect 479 365 483 369
rect 485 365 489 369
rect 491 365 495 369
rect 497 365 501 369
rect 503 365 507 369
rect 509 365 513 369
rect 515 365 519 369
rect 521 365 525 369
rect 527 365 531 369
rect 533 365 537 369
rect 539 365 543 369
rect 545 365 549 369
rect 551 365 555 369
rect 557 365 561 369
rect 563 365 567 369
rect 569 365 573 369
rect 575 365 579 369
rect 581 365 585 369
rect 587 365 591 369
rect 617 365 621 369
rect 623 365 627 369
rect 629 365 633 369
rect 635 365 639 369
rect 641 365 645 369
rect 647 365 651 369
rect 653 365 657 369
rect 659 365 663 369
rect 665 365 669 369
rect 671 365 675 369
rect 677 365 681 369
rect 683 365 687 369
rect 689 365 693 369
rect 695 365 699 369
rect 701 365 705 369
rect 707 365 711 369
rect 713 365 717 369
rect 719 365 723 369
rect 725 365 729 369
rect 731 365 735 369
rect 737 365 741 369
rect 743 365 747 369
rect 749 365 753 369
rect 755 365 759 369
rect 761 365 765 369
rect 767 365 771 369
rect 773 365 777 369
rect 779 365 783 369
rect 785 365 789 369
rect 791 365 795 369
rect 797 365 801 369
rect 803 365 807 369
rect 809 365 813 369
rect 815 365 819 369
rect 821 365 825 369
rect 827 365 831 369
rect 833 365 837 369
rect 839 365 843 369
rect 845 365 849 369
rect 851 365 855 369
rect 857 365 861 369
rect 863 365 867 369
rect 869 365 873 369
rect 875 365 879 369
rect 881 365 885 369
rect 887 365 891 369
rect 893 365 897 369
rect 899 365 903 369
rect 905 365 909 369
rect 911 365 915 369
rect 917 365 921 369
rect 923 365 927 369
rect 929 365 933 369
rect 935 365 939 369
rect 941 365 945 369
rect 947 365 951 369
rect 953 365 957 369
rect 959 365 963 369
rect 965 365 969 369
rect 971 365 975 369
rect 977 365 981 369
rect 983 365 987 369
rect 989 365 993 369
rect 995 365 999 369
rect 1001 365 1005 369
rect 1007 365 1011 369
rect 1013 365 1017 369
rect 1019 365 1023 369
rect 1025 365 1029 369
rect 1031 365 1035 369
rect 1037 365 1041 369
rect 1043 365 1047 369
rect 1049 365 1053 369
rect 1055 365 1059 369
rect 1061 365 1065 369
rect 1091 365 1095 369
rect 1097 365 1101 369
rect 1103 365 1107 369
rect 1109 365 1113 369
rect 1115 365 1119 369
rect 1121 365 1125 369
rect 1127 365 1131 369
rect 1133 365 1137 369
rect 1139 365 1143 369
rect 1145 365 1149 369
rect 1151 365 1155 369
rect 1157 365 1161 369
rect 1163 365 1167 369
rect 1169 365 1173 369
rect 1175 365 1179 369
rect 1181 365 1185 369
rect 1187 365 1191 369
rect 1193 365 1197 369
rect 1199 365 1203 369
rect 1205 365 1209 369
rect 1211 365 1215 369
rect 1217 365 1221 369
rect 1223 365 1227 369
rect 1229 365 1233 369
rect 1235 365 1239 369
rect 1241 365 1245 369
rect 1247 365 1251 369
rect 1253 365 1257 369
rect 1259 365 1263 369
rect 1265 365 1269 369
rect 1271 365 1275 369
rect 1277 365 1281 369
rect 1283 365 1287 369
rect 1289 365 1293 369
rect 1295 365 1299 369
rect 1301 365 1305 369
rect 1307 365 1311 369
rect 1313 365 1317 369
rect 1319 365 1323 369
rect 1325 365 1329 369
rect 1331 365 1335 369
rect 1337 365 1341 369
rect 1343 365 1347 369
rect 1349 365 1353 369
rect 1355 365 1359 369
rect 1361 365 1365 369
rect 1367 365 1371 369
rect 1373 365 1377 369
rect 1379 365 1383 369
rect 1385 365 1389 369
rect 1391 365 1395 369
rect 1397 365 1401 369
rect 1403 365 1407 369
rect 1409 365 1413 369
rect 1415 365 1419 369
rect 1421 365 1425 369
rect 1427 365 1431 369
rect 1433 365 1437 369
rect 1439 365 1443 369
rect 1445 365 1449 369
rect 1451 365 1455 369
rect 1457 365 1461 369
rect 1463 365 1467 369
rect 1469 365 1473 369
rect 1475 365 1479 369
rect 1481 365 1485 369
rect 1487 365 1491 369
rect 1493 365 1497 369
rect 1499 365 1503 369
rect 1505 365 1509 369
rect 1511 365 1515 369
rect 1517 365 1521 369
rect 1523 365 1527 369
rect 1529 365 1533 369
rect 1535 365 1539 369
rect 1565 365 1569 369
rect 1571 365 1575 369
rect 1577 365 1581 369
rect 1583 365 1587 369
rect 1589 365 1593 369
rect 1595 365 1599 369
rect 1601 365 1605 369
rect 1607 365 1611 369
rect 1613 365 1617 369
rect 1619 365 1623 369
rect 1625 365 1629 369
rect 1631 365 1635 369
rect 1637 365 1641 369
rect 1643 365 1647 369
rect 1649 365 1653 369
rect 1655 365 1659 369
rect 1661 365 1665 369
rect 1667 365 1671 369
rect 1673 365 1677 369
rect 1679 365 1683 369
rect 1685 365 1689 369
rect 1691 365 1695 369
rect 1697 365 1701 369
rect 1703 365 1707 369
rect 1709 365 1713 369
rect 1715 365 1719 369
rect 1721 365 1725 369
rect 1727 365 1731 369
rect 1733 365 1737 369
rect 1739 365 1743 369
rect 1745 365 1749 369
rect 1751 365 1755 369
rect 1757 365 1761 369
rect 1763 365 1767 369
rect 1769 365 1773 369
rect 1775 365 1779 369
rect 1781 365 1785 369
rect 1787 365 1791 369
rect 1793 365 1797 369
rect 1799 365 1803 369
rect 1805 365 1809 369
rect 1811 365 1815 369
rect 1817 365 1821 369
rect 1823 365 1827 369
rect 1829 365 1833 369
rect 1835 365 1839 369
rect 1841 365 1845 369
rect 1847 365 1851 369
rect 1853 365 1857 369
rect 1859 365 1863 369
rect 1865 365 1869 369
rect 1871 365 1875 369
rect 1877 365 1881 369
rect 1883 365 1887 369
rect 1889 365 1893 369
rect 1895 365 1899 369
rect 1901 365 1905 369
rect 1907 365 1911 369
rect 1913 365 1917 369
rect 1919 365 1923 369
rect 1925 365 1929 369
rect 1931 365 1935 369
rect 1937 365 1941 369
rect 1943 365 1947 369
rect 1949 365 1953 369
rect 1955 365 1959 369
rect 1961 365 1965 369
rect 1967 365 1971 369
rect 1973 365 1977 369
rect 1979 365 1983 369
rect 1985 365 1989 369
rect 1991 365 1995 369
rect 1997 365 2001 369
rect 2003 365 2007 369
rect 2009 365 2013 369
rect 2039 365 2043 369
rect 2045 365 2049 369
rect 2051 365 2055 369
rect 2057 365 2061 369
rect 2063 365 2067 369
rect 2069 365 2073 369
rect 2075 365 2079 369
rect 2081 365 2085 369
rect 2087 365 2091 369
rect 2093 365 2097 369
rect 2099 365 2103 369
rect 2105 365 2109 369
rect 2111 365 2115 369
rect 2117 365 2121 369
rect 2123 365 2127 369
rect 2129 365 2133 369
rect 2135 365 2139 369
rect 2141 365 2145 369
rect 2147 365 2151 369
rect 2153 365 2157 369
rect 2159 365 2163 369
rect 2165 365 2169 369
rect 2171 365 2175 369
rect 2177 365 2181 369
rect 2183 365 2187 369
rect 2189 365 2193 369
rect 2195 365 2199 369
rect 2201 365 2205 369
rect 2207 365 2211 369
rect 2213 365 2217 369
rect 2219 365 2223 369
rect 2225 365 2229 369
rect 2231 365 2235 369
rect 2237 365 2241 369
rect 2243 365 2247 369
rect 2249 365 2253 369
rect 2255 365 2259 369
rect 2261 365 2265 369
rect 2267 365 2271 369
rect 2273 365 2277 369
rect 2279 365 2283 369
rect 2285 365 2289 369
rect 2291 365 2295 369
rect 2297 365 2301 369
rect 2303 365 2307 369
rect 2309 365 2313 369
rect 2315 365 2319 369
rect 2321 365 2325 369
rect 2327 365 2331 369
rect 2333 365 2337 369
rect 2339 365 2343 369
rect 2345 365 2349 369
rect 2351 365 2355 369
rect 2357 365 2361 369
rect 2363 365 2367 369
rect 2369 365 2373 369
rect 2375 365 2379 369
rect 2381 365 2385 369
rect 2387 365 2391 369
rect 2393 365 2397 369
rect 2399 365 2403 369
rect 2405 365 2409 369
rect 2411 365 2415 369
rect 2417 365 2421 369
rect 2423 365 2427 369
rect 2429 365 2433 369
rect 2435 365 2439 369
rect 2441 365 2445 369
rect 2447 365 2451 369
rect 2453 365 2457 369
rect 2459 365 2463 369
rect 2465 365 2469 369
rect 2471 365 2475 369
rect 2477 365 2481 369
rect 2483 365 2487 369
rect 2513 365 2517 369
rect 2519 365 2523 369
rect 2525 365 2529 369
rect 2531 365 2535 369
rect 2537 365 2541 369
rect 2543 365 2547 369
rect 2549 365 2553 369
rect 2555 365 2559 369
rect 2561 365 2565 369
rect 2567 365 2571 369
rect 2573 365 2577 369
rect 2579 365 2583 369
rect 2585 365 2589 369
rect 2591 365 2595 369
rect 2597 365 2601 369
rect 2603 365 2607 369
rect 2609 365 2613 369
rect 2615 365 2619 369
rect 2621 365 2625 369
rect 2627 365 2631 369
rect 2633 365 2637 369
rect 2639 365 2643 369
rect 2645 365 2649 369
rect 2651 365 2655 369
rect 2657 365 2661 369
rect 2663 365 2667 369
rect 2669 365 2673 369
rect 2675 365 2679 369
rect 2681 365 2685 369
rect 2687 365 2691 369
rect 2693 365 2697 369
rect 2699 365 2703 369
rect 2705 365 2709 369
rect 2711 365 2715 369
rect 2717 365 2721 369
rect 2723 365 2727 369
rect 2729 365 2733 369
rect 2735 365 2739 369
rect 2741 365 2745 369
rect 2747 365 2751 369
rect 2753 365 2757 369
rect 2759 365 2763 369
rect 2765 365 2769 369
rect 2771 365 2775 369
rect 2777 365 2781 369
rect 2783 365 2787 369
rect 2789 365 2793 369
rect 2795 365 2799 369
rect 2801 365 2805 369
rect 2807 365 2811 369
rect 2813 365 2817 369
rect 2819 365 2823 369
rect 2825 365 2829 369
rect 2831 365 2835 369
rect 2837 365 2841 369
rect 2843 365 2847 369
rect 2849 365 2853 369
rect 2855 365 2859 369
rect 2861 365 2865 369
rect 2867 365 2871 369
rect 2873 365 2877 369
rect 2879 365 2883 369
rect 2885 365 2889 369
rect 2891 365 2895 369
rect 2897 365 2901 369
rect 2903 365 2907 369
rect 2909 365 2913 369
rect 2915 365 2919 369
rect 2921 365 2925 369
rect 2927 365 2931 369
rect 2933 365 2937 369
rect 2939 365 2943 369
rect 2945 365 2949 369
rect 2951 365 2955 369
rect 2957 365 2961 369
rect 2987 365 2991 369
rect 2993 365 2997 369
rect 2999 365 3003 369
rect 3005 365 3009 369
rect 3011 365 3015 369
rect 3017 365 3021 369
rect 3023 365 3027 369
rect 3029 365 3033 369
rect 3035 365 3039 369
rect 3041 365 3045 369
rect 3047 365 3051 369
rect 3053 365 3057 369
rect 3059 365 3063 369
rect 3065 365 3069 369
rect 3071 365 3075 369
rect 3077 365 3081 369
rect 3083 365 3087 369
rect 3089 365 3093 369
rect 3095 365 3099 369
rect 3101 365 3105 369
rect 3107 365 3111 369
rect 3113 365 3117 369
rect 3119 365 3123 369
rect 3125 365 3129 369
rect 3131 365 3135 369
rect 3137 365 3141 369
rect 3143 365 3147 369
rect 3149 365 3153 369
rect 3155 365 3159 369
rect 3161 365 3165 369
rect 3167 365 3171 369
rect 3173 365 3177 369
rect 3179 365 3183 369
rect 3185 365 3189 369
rect 3191 365 3195 369
rect 3197 365 3201 369
rect 3203 365 3207 369
rect 3209 365 3213 369
rect 3215 365 3219 369
rect 3221 365 3225 369
rect 3227 365 3231 369
rect 3233 365 3237 369
rect 3239 365 3243 369
rect 3245 365 3249 369
rect 3251 365 3255 369
rect 3257 365 3261 369
rect 3263 365 3267 369
rect 3269 365 3273 369
rect 3275 365 3279 369
rect 3281 365 3285 369
rect 3287 365 3291 369
rect 3293 365 3297 369
rect 3299 365 3303 369
rect 3305 365 3309 369
rect 3311 365 3315 369
rect 3317 365 3321 369
rect 3323 365 3327 369
rect 3329 365 3333 369
rect 3335 365 3339 369
rect 3341 365 3345 369
rect 3347 365 3351 369
rect 3353 365 3357 369
rect 3359 365 3363 369
rect 3365 365 3369 369
rect 3371 365 3375 369
rect 3377 365 3381 369
rect 3383 365 3387 369
rect 3389 365 3393 369
rect 3395 365 3399 369
rect 3401 365 3405 369
rect 3407 365 3411 369
rect 3413 365 3417 369
rect 3419 365 3423 369
rect 3425 365 3429 369
rect 3431 365 3435 369
rect 3461 365 3465 369
rect 3467 365 3471 369
rect 3473 365 3477 369
rect 3479 365 3483 369
rect 3485 365 3489 369
rect 3491 365 3495 369
rect 3497 365 3501 369
rect 3503 365 3507 369
rect 3509 365 3513 369
rect 3515 365 3519 369
rect 3521 365 3525 369
rect 3527 365 3531 369
rect 3533 365 3537 369
rect 3539 365 3543 369
rect 3545 365 3549 369
rect 3551 365 3555 369
rect 3557 365 3561 369
rect 3563 365 3567 369
rect 3569 365 3573 369
rect 3575 365 3579 369
rect 3581 365 3585 369
rect 3587 365 3591 369
rect 3593 365 3597 369
rect 3599 365 3603 369
rect 3605 365 3609 369
rect 3611 365 3615 369
rect 3617 365 3621 369
rect 3623 365 3627 369
rect 3629 365 3633 369
rect 3635 365 3639 369
rect 3641 365 3645 369
rect 3647 365 3651 369
rect 3653 365 3657 369
rect 3659 365 3663 369
rect 3665 365 3669 369
rect 3671 365 3675 369
rect 3677 365 3681 369
rect 3683 365 3687 369
rect 3689 365 3693 369
rect 3695 365 3699 369
rect 3701 365 3705 369
rect 3707 365 3711 369
rect 3713 365 3717 369
rect 3719 365 3723 369
rect 3725 365 3729 369
rect 3731 365 3735 369
rect 3737 365 3741 369
rect 3743 365 3747 369
rect 3749 365 3753 369
rect 3755 365 3759 369
rect 3761 365 3765 369
rect 3767 365 3771 369
rect 3773 365 3777 369
rect 3779 365 3783 369
rect 3785 365 3789 369
rect 3791 365 3795 369
rect 3797 365 3801 369
rect 3803 365 3807 369
rect 3809 365 3813 369
rect 3815 365 3819 369
rect 3821 365 3825 369
rect 3827 365 3831 369
rect 3833 365 3837 369
rect 3839 365 3843 369
rect 3845 365 3849 369
rect 3851 365 3855 369
rect 3857 365 3861 369
rect 3863 365 3867 369
rect 3869 365 3873 369
rect 3875 365 3879 369
rect 3881 365 3885 369
rect 3887 365 3891 369
rect 3893 365 3897 369
rect 3899 365 3903 369
rect 3905 365 3909 369
rect 3935 365 3939 369
rect 3941 365 3945 369
rect 3947 365 3951 369
rect 3953 365 3957 369
rect 3959 365 3963 369
rect 3965 365 3969 369
rect 3971 365 3975 369
rect 3977 365 3981 369
rect 3983 365 3987 369
rect 3989 365 3993 369
rect 3995 365 3999 369
rect 4001 365 4005 369
rect 4007 365 4011 369
rect 4013 365 4017 369
rect 4019 365 4023 369
rect 4025 365 4029 369
rect 4031 365 4035 369
rect 4037 365 4041 369
rect 4043 365 4047 369
rect 4049 365 4053 369
rect 4055 365 4059 369
rect 4061 365 4065 369
rect 4067 365 4071 369
rect 4073 365 4077 369
rect 4079 365 4083 369
rect 4085 365 4089 369
rect 4091 365 4095 369
rect 4097 365 4101 369
rect 4103 365 4107 369
rect 4109 365 4113 369
rect 4115 365 4119 369
rect 4121 365 4125 369
rect 4127 365 4131 369
rect 4133 365 4137 369
rect 4139 365 4143 369
rect 4145 365 4149 369
rect 4151 365 4155 369
rect 4157 365 4161 369
rect 4163 365 4167 369
rect 4169 365 4173 369
rect 4175 365 4179 369
rect 4181 365 4185 369
rect 4187 365 4191 369
rect 4193 365 4197 369
rect 4199 365 4203 369
rect 4205 365 4209 369
rect 4211 365 4215 369
rect 4217 365 4221 369
rect 4223 365 4227 369
rect 4229 365 4233 369
rect 4235 365 4239 369
rect 4241 365 4245 369
rect 4247 365 4251 369
rect 4253 365 4257 369
rect 4259 365 4263 369
rect 4265 365 4269 369
rect 4271 365 4275 369
rect 4277 365 4281 369
rect 4283 365 4287 369
rect 4289 365 4293 369
rect 4295 365 4299 369
rect 4301 365 4305 369
rect 4307 365 4311 369
rect 4313 365 4317 369
rect 4319 365 4323 369
rect 4325 365 4329 369
rect 4331 365 4335 369
rect 4337 365 4341 369
rect 4343 365 4347 369
rect 4349 365 4353 369
rect 4355 365 4359 369
rect 4361 365 4365 369
rect 4367 365 4371 369
rect 4373 365 4377 369
rect 4379 365 4383 369
rect 4409 365 4413 369
rect 4415 365 4419 369
rect 4421 365 4425 369
rect 4427 365 4431 369
rect 4433 365 4437 369
rect 4439 365 4443 369
rect 4445 365 4449 369
rect 4451 365 4455 369
rect 4457 365 4461 369
rect 4463 365 4467 369
rect 4469 365 4473 369
rect 4475 365 4479 369
rect 4481 365 4485 369
rect 4487 365 4491 369
rect 4493 365 4497 369
rect 4499 365 4503 369
rect 4505 365 4509 369
rect 4511 365 4515 369
rect 4517 365 4521 369
rect 4523 365 4527 369
rect 4529 365 4533 369
rect 4535 365 4539 369
rect 4541 365 4545 369
rect 4547 365 4551 369
rect 4553 365 4557 369
rect 4559 365 4563 369
rect 4565 365 4569 369
rect 4571 365 4575 369
rect 4577 365 4581 369
rect 4583 365 4587 369
rect 4589 365 4593 369
rect 4595 365 4599 369
rect 4601 365 4605 369
rect 4607 365 4611 369
rect 4613 365 4617 369
rect 4619 365 4623 369
rect 4625 365 4629 369
rect 4631 365 4635 369
rect 4637 365 4641 369
rect 4643 365 4647 369
rect 4649 365 4653 369
rect 4655 365 4659 369
rect 4661 365 4665 369
rect 4667 365 4671 369
rect 4673 365 4677 369
rect 4679 365 4683 369
rect 4685 365 4689 369
rect 4691 365 4695 369
rect 4697 365 4701 369
rect 4703 365 4707 369
rect 4709 365 4713 369
rect 4715 365 4719 369
rect 4721 365 4725 369
rect 4727 365 4731 369
rect 4733 365 4737 369
rect 4739 365 4743 369
rect 4745 365 4749 369
rect 4751 365 4755 369
rect 4757 365 4761 369
rect 4763 365 4767 369
rect 4769 365 4773 369
rect 4775 365 4779 369
rect 4781 365 4785 369
rect 4787 365 4791 369
rect 4793 365 4797 369
rect 4799 365 4803 369
rect 4805 365 4809 369
rect 4811 365 4815 369
rect 4817 365 4821 369
rect 4823 365 4827 369
rect 4829 365 4833 369
rect 4835 365 4839 369
rect 4841 365 4845 369
rect 4847 365 4851 369
rect 4853 365 4857 369
rect 4859 365 4863 369
rect 4865 365 4869 369
rect 4871 365 4875 369
rect 4877 365 4881 369
rect 4883 365 4887 369
rect 4889 365 4893 369
rect 4895 365 4899 369
rect 4901 365 4905 369
rect 4907 365 4911 369
rect 4913 365 4917 369
rect 4919 365 4923 369
rect 4925 365 4929 369
rect 4931 365 4935 369
rect 4937 365 4941 369
rect 4943 365 4947 369
rect 4949 365 4953 369
rect 4955 365 4959 369
rect 4961 365 4965 369
rect 4967 365 4971 369
rect 4973 365 4977 369
rect 4979 365 4983 369
rect 4985 365 4989 369
rect 4991 365 4995 369
rect 365 359 369 363
rect 365 353 369 357
rect 365 347 369 351
rect 365 341 369 345
rect 365 335 369 339
rect 365 329 369 333
rect 365 323 369 327
rect 365 317 369 321
rect 365 311 369 315
rect 365 305 369 309
rect 365 299 369 303
rect 365 293 369 297
rect 365 287 369 291
rect 365 281 369 285
rect 365 275 369 279
rect 365 269 369 273
rect 365 263 369 267
rect 365 257 369 261
rect 365 251 369 255
rect 365 245 369 249
rect 365 239 369 243
rect 365 233 369 237
rect 365 227 369 231
rect 365 221 369 225
rect 365 215 369 219
rect 365 209 369 213
rect 365 203 369 207
rect 365 197 369 201
rect 365 191 369 195
rect 365 185 369 189
rect 365 179 369 183
rect 365 173 369 177
rect 365 167 369 171
rect 365 161 369 165
rect 365 155 369 159
rect 365 149 369 153
rect 365 143 369 147
rect 365 137 369 141
rect 365 131 369 135
rect 365 125 369 129
rect 365 119 369 123
rect 365 113 369 117
rect 365 107 369 111
rect 365 101 369 105
rect 365 95 369 99
rect 365 89 369 93
rect 365 83 369 87
rect 365 77 369 81
rect 365 71 369 75
rect 365 65 369 69
rect 365 59 369 63
rect 365 53 369 57
rect 365 47 369 51
rect 365 41 369 45
rect 365 35 369 39
rect 365 29 369 33
rect 365 23 369 27
rect 365 17 369 21
rect 365 11 369 15
rect 365 5 369 9
rect 839 359 843 363
rect 839 353 843 357
rect 839 347 843 351
rect 839 341 843 345
rect 839 335 843 339
rect 839 329 843 333
rect 839 323 843 327
rect 839 317 843 321
rect 839 311 843 315
rect 839 305 843 309
rect 839 299 843 303
rect 839 293 843 297
rect 839 287 843 291
rect 839 281 843 285
rect 839 275 843 279
rect 839 269 843 273
rect 839 263 843 267
rect 839 257 843 261
rect 839 251 843 255
rect 839 245 843 249
rect 839 239 843 243
rect 839 233 843 237
rect 839 227 843 231
rect 839 221 843 225
rect 839 215 843 219
rect 839 209 843 213
rect 839 203 843 207
rect 839 197 843 201
rect 839 191 843 195
rect 839 185 843 189
rect 839 179 843 183
rect 839 173 843 177
rect 839 167 843 171
rect 839 161 843 165
rect 839 155 843 159
rect 839 149 843 153
rect 839 143 843 147
rect 839 137 843 141
rect 839 131 843 135
rect 839 125 843 129
rect 839 119 843 123
rect 839 113 843 117
rect 839 107 843 111
rect 839 101 843 105
rect 839 95 843 99
rect 839 89 843 93
rect 839 83 843 87
rect 839 77 843 81
rect 839 71 843 75
rect 839 65 843 69
rect 839 59 843 63
rect 839 53 843 57
rect 839 47 843 51
rect 839 41 843 45
rect 839 35 843 39
rect 839 29 843 33
rect 839 23 843 27
rect 839 17 843 21
rect 839 11 843 15
rect 839 5 843 9
rect 1313 359 1317 363
rect 1313 353 1317 357
rect 1313 347 1317 351
rect 1313 341 1317 345
rect 1313 335 1317 339
rect 1313 329 1317 333
rect 1313 323 1317 327
rect 1313 317 1317 321
rect 1313 311 1317 315
rect 1313 305 1317 309
rect 1313 299 1317 303
rect 1313 293 1317 297
rect 1313 287 1317 291
rect 1313 281 1317 285
rect 1313 275 1317 279
rect 1313 269 1317 273
rect 1313 263 1317 267
rect 1313 257 1317 261
rect 1313 251 1317 255
rect 1313 245 1317 249
rect 1313 239 1317 243
rect 1313 233 1317 237
rect 1313 227 1317 231
rect 1313 221 1317 225
rect 1313 215 1317 219
rect 1313 209 1317 213
rect 1313 203 1317 207
rect 1313 197 1317 201
rect 1313 191 1317 195
rect 1313 185 1317 189
rect 1313 179 1317 183
rect 1313 173 1317 177
rect 1313 167 1317 171
rect 1313 161 1317 165
rect 1313 155 1317 159
rect 1313 149 1317 153
rect 1313 143 1317 147
rect 1313 137 1317 141
rect 1313 131 1317 135
rect 1313 125 1317 129
rect 1313 119 1317 123
rect 1313 113 1317 117
rect 1313 107 1317 111
rect 1313 101 1317 105
rect 1313 95 1317 99
rect 1313 89 1317 93
rect 1313 83 1317 87
rect 1313 77 1317 81
rect 1313 71 1317 75
rect 1313 65 1317 69
rect 1313 59 1317 63
rect 1313 53 1317 57
rect 1313 47 1317 51
rect 1313 41 1317 45
rect 1313 35 1317 39
rect 1313 29 1317 33
rect 1313 23 1317 27
rect 1313 17 1317 21
rect 1313 11 1317 15
rect 1313 5 1317 9
rect 1787 359 1791 363
rect 1787 353 1791 357
rect 1787 347 1791 351
rect 1787 341 1791 345
rect 1787 335 1791 339
rect 1787 329 1791 333
rect 1787 323 1791 327
rect 1787 317 1791 321
rect 1787 311 1791 315
rect 1787 305 1791 309
rect 1787 299 1791 303
rect 1787 293 1791 297
rect 1787 287 1791 291
rect 1787 281 1791 285
rect 1787 275 1791 279
rect 1787 269 1791 273
rect 1787 263 1791 267
rect 1787 257 1791 261
rect 1787 251 1791 255
rect 1787 245 1791 249
rect 1787 239 1791 243
rect 1787 233 1791 237
rect 1787 227 1791 231
rect 1787 221 1791 225
rect 1787 215 1791 219
rect 1787 209 1791 213
rect 1787 203 1791 207
rect 1787 197 1791 201
rect 1787 191 1791 195
rect 1787 185 1791 189
rect 1787 179 1791 183
rect 1787 173 1791 177
rect 1787 167 1791 171
rect 1787 161 1791 165
rect 1787 155 1791 159
rect 1787 149 1791 153
rect 1787 143 1791 147
rect 1787 137 1791 141
rect 1787 131 1791 135
rect 1787 125 1791 129
rect 1787 119 1791 123
rect 1787 113 1791 117
rect 1787 107 1791 111
rect 1787 101 1791 105
rect 1787 95 1791 99
rect 1787 89 1791 93
rect 1787 83 1791 87
rect 1787 77 1791 81
rect 1787 71 1791 75
rect 1787 65 1791 69
rect 1787 59 1791 63
rect 1787 53 1791 57
rect 1787 47 1791 51
rect 1787 41 1791 45
rect 1787 35 1791 39
rect 1787 29 1791 33
rect 1787 23 1791 27
rect 1787 17 1791 21
rect 1787 11 1791 15
rect 1787 5 1791 9
rect 2261 359 2265 363
rect 2261 353 2265 357
rect 2261 347 2265 351
rect 2261 341 2265 345
rect 2261 335 2265 339
rect 2261 329 2265 333
rect 2261 323 2265 327
rect 2261 317 2265 321
rect 2261 311 2265 315
rect 2261 305 2265 309
rect 2261 299 2265 303
rect 2261 293 2265 297
rect 2261 287 2265 291
rect 2261 281 2265 285
rect 2261 275 2265 279
rect 2261 269 2265 273
rect 2261 263 2265 267
rect 2261 257 2265 261
rect 2261 251 2265 255
rect 2261 245 2265 249
rect 2261 239 2265 243
rect 2261 233 2265 237
rect 2261 227 2265 231
rect 2261 221 2265 225
rect 2261 215 2265 219
rect 2261 209 2265 213
rect 2261 203 2265 207
rect 2261 197 2265 201
rect 2261 191 2265 195
rect 2261 185 2265 189
rect 2261 179 2265 183
rect 2261 173 2265 177
rect 2261 167 2265 171
rect 2261 161 2265 165
rect 2261 155 2265 159
rect 2261 149 2265 153
rect 2261 143 2265 147
rect 2261 137 2265 141
rect 2261 131 2265 135
rect 2261 125 2265 129
rect 2261 119 2265 123
rect 2261 113 2265 117
rect 2261 107 2265 111
rect 2261 101 2265 105
rect 2261 95 2265 99
rect 2261 89 2265 93
rect 2261 83 2265 87
rect 2261 77 2265 81
rect 2261 71 2265 75
rect 2261 65 2265 69
rect 2261 59 2265 63
rect 2261 53 2265 57
rect 2261 47 2265 51
rect 2261 41 2265 45
rect 2261 35 2265 39
rect 2261 29 2265 33
rect 2261 23 2265 27
rect 2261 17 2265 21
rect 2261 11 2265 15
rect 2261 5 2265 9
rect 2735 359 2739 363
rect 2735 353 2739 357
rect 2735 347 2739 351
rect 2735 341 2739 345
rect 2735 335 2739 339
rect 2735 329 2739 333
rect 2735 323 2739 327
rect 2735 317 2739 321
rect 2735 311 2739 315
rect 2735 305 2739 309
rect 2735 299 2739 303
rect 2735 293 2739 297
rect 2735 287 2739 291
rect 2735 281 2739 285
rect 2735 275 2739 279
rect 2735 269 2739 273
rect 2735 263 2739 267
rect 2735 257 2739 261
rect 2735 251 2739 255
rect 2735 245 2739 249
rect 2735 239 2739 243
rect 2735 233 2739 237
rect 2735 227 2739 231
rect 2735 221 2739 225
rect 2735 215 2739 219
rect 2735 209 2739 213
rect 2735 203 2739 207
rect 2735 197 2739 201
rect 2735 191 2739 195
rect 2735 185 2739 189
rect 2735 179 2739 183
rect 2735 173 2739 177
rect 2735 167 2739 171
rect 2735 161 2739 165
rect 2735 155 2739 159
rect 2735 149 2739 153
rect 2735 143 2739 147
rect 2735 137 2739 141
rect 2735 131 2739 135
rect 2735 125 2739 129
rect 2735 119 2739 123
rect 2735 113 2739 117
rect 2735 107 2739 111
rect 2735 101 2739 105
rect 2735 95 2739 99
rect 2735 89 2739 93
rect 2735 83 2739 87
rect 2735 77 2739 81
rect 2735 71 2739 75
rect 2735 65 2739 69
rect 2735 59 2739 63
rect 2735 53 2739 57
rect 2735 47 2739 51
rect 2735 41 2739 45
rect 2735 35 2739 39
rect 2735 29 2739 33
rect 2735 23 2739 27
rect 2735 17 2739 21
rect 2735 11 2739 15
rect 2735 5 2739 9
rect 3209 359 3213 363
rect 3209 353 3213 357
rect 3209 347 3213 351
rect 3209 341 3213 345
rect 3209 335 3213 339
rect 3209 329 3213 333
rect 3209 323 3213 327
rect 3209 317 3213 321
rect 3209 311 3213 315
rect 3209 305 3213 309
rect 3209 299 3213 303
rect 3209 293 3213 297
rect 3209 287 3213 291
rect 3209 281 3213 285
rect 3209 275 3213 279
rect 3209 269 3213 273
rect 3209 263 3213 267
rect 3209 257 3213 261
rect 3209 251 3213 255
rect 3209 245 3213 249
rect 3209 239 3213 243
rect 3209 233 3213 237
rect 3209 227 3213 231
rect 3209 221 3213 225
rect 3209 215 3213 219
rect 3209 209 3213 213
rect 3209 203 3213 207
rect 3209 197 3213 201
rect 3209 191 3213 195
rect 3209 185 3213 189
rect 3209 179 3213 183
rect 3209 173 3213 177
rect 3209 167 3213 171
rect 3209 161 3213 165
rect 3209 155 3213 159
rect 3209 149 3213 153
rect 3209 143 3213 147
rect 3209 137 3213 141
rect 3209 131 3213 135
rect 3209 125 3213 129
rect 3209 119 3213 123
rect 3209 113 3213 117
rect 3209 107 3213 111
rect 3209 101 3213 105
rect 3209 95 3213 99
rect 3209 89 3213 93
rect 3209 83 3213 87
rect 3209 77 3213 81
rect 3209 71 3213 75
rect 3209 65 3213 69
rect 3209 59 3213 63
rect 3209 53 3213 57
rect 3209 47 3213 51
rect 3209 41 3213 45
rect 3209 35 3213 39
rect 3209 29 3213 33
rect 3209 23 3213 27
rect 3209 17 3213 21
rect 3209 11 3213 15
rect 3209 5 3213 9
rect 3683 359 3687 363
rect 3683 353 3687 357
rect 3683 347 3687 351
rect 3683 341 3687 345
rect 3683 335 3687 339
rect 3683 329 3687 333
rect 3683 323 3687 327
rect 3683 317 3687 321
rect 3683 311 3687 315
rect 3683 305 3687 309
rect 3683 299 3687 303
rect 3683 293 3687 297
rect 3683 287 3687 291
rect 3683 281 3687 285
rect 3683 275 3687 279
rect 3683 269 3687 273
rect 3683 263 3687 267
rect 3683 257 3687 261
rect 3683 251 3687 255
rect 3683 245 3687 249
rect 3683 239 3687 243
rect 3683 233 3687 237
rect 3683 227 3687 231
rect 3683 221 3687 225
rect 3683 215 3687 219
rect 3683 209 3687 213
rect 3683 203 3687 207
rect 3683 197 3687 201
rect 3683 191 3687 195
rect 3683 185 3687 189
rect 3683 179 3687 183
rect 3683 173 3687 177
rect 3683 167 3687 171
rect 3683 161 3687 165
rect 3683 155 3687 159
rect 3683 149 3687 153
rect 3683 143 3687 147
rect 3683 137 3687 141
rect 3683 131 3687 135
rect 3683 125 3687 129
rect 3683 119 3687 123
rect 3683 113 3687 117
rect 3683 107 3687 111
rect 3683 101 3687 105
rect 3683 95 3687 99
rect 3683 89 3687 93
rect 3683 83 3687 87
rect 3683 77 3687 81
rect 3683 71 3687 75
rect 3683 65 3687 69
rect 3683 59 3687 63
rect 3683 53 3687 57
rect 3683 47 3687 51
rect 3683 41 3687 45
rect 3683 35 3687 39
rect 3683 29 3687 33
rect 3683 23 3687 27
rect 3683 17 3687 21
rect 3683 11 3687 15
rect 3683 5 3687 9
rect 4157 359 4161 363
rect 4157 353 4161 357
rect 4157 347 4161 351
rect 4157 341 4161 345
rect 4157 335 4161 339
rect 4157 329 4161 333
rect 4157 323 4161 327
rect 4157 317 4161 321
rect 4157 311 4161 315
rect 4157 305 4161 309
rect 4157 299 4161 303
rect 4157 293 4161 297
rect 4157 287 4161 291
rect 4157 281 4161 285
rect 4157 275 4161 279
rect 4157 269 4161 273
rect 4157 263 4161 267
rect 4157 257 4161 261
rect 4157 251 4161 255
rect 4157 245 4161 249
rect 4157 239 4161 243
rect 4157 233 4161 237
rect 4157 227 4161 231
rect 4157 221 4161 225
rect 4157 215 4161 219
rect 4157 209 4161 213
rect 4157 203 4161 207
rect 4157 197 4161 201
rect 4157 191 4161 195
rect 4157 185 4161 189
rect 4157 179 4161 183
rect 4157 173 4161 177
rect 4157 167 4161 171
rect 4157 161 4161 165
rect 4157 155 4161 159
rect 4157 149 4161 153
rect 4157 143 4161 147
rect 4157 137 4161 141
rect 4157 131 4161 135
rect 4157 125 4161 129
rect 4157 119 4161 123
rect 4157 113 4161 117
rect 4157 107 4161 111
rect 4157 101 4161 105
rect 4157 95 4161 99
rect 4157 89 4161 93
rect 4157 83 4161 87
rect 4157 77 4161 81
rect 4157 71 4161 75
rect 4157 65 4161 69
rect 4157 59 4161 63
rect 4157 53 4161 57
rect 4157 47 4161 51
rect 4157 41 4161 45
rect 4157 35 4161 39
rect 4157 29 4161 33
rect 4157 23 4161 27
rect 4157 17 4161 21
rect 4157 11 4161 15
rect 4157 5 4161 9
rect 4631 359 4635 363
rect 4631 353 4635 357
rect 4631 347 4635 351
rect 4631 341 4635 345
rect 4631 335 4635 339
rect 4631 329 4635 333
rect 4631 323 4635 327
rect 4631 317 4635 321
rect 4631 311 4635 315
rect 4631 305 4635 309
rect 4631 299 4635 303
rect 4631 293 4635 297
rect 4631 287 4635 291
rect 4631 281 4635 285
rect 4631 275 4635 279
rect 4631 269 4635 273
rect 4631 263 4635 267
rect 4631 257 4635 261
rect 4631 251 4635 255
rect 4631 245 4635 249
rect 4631 239 4635 243
rect 4631 233 4635 237
rect 4631 227 4635 231
rect 4631 221 4635 225
rect 4631 215 4635 219
rect 4631 209 4635 213
rect 4631 203 4635 207
rect 4631 197 4635 201
rect 4631 191 4635 195
rect 4631 185 4635 189
rect 4631 179 4635 183
rect 4631 173 4635 177
rect 4631 167 4635 171
rect 4631 161 4635 165
rect 4631 155 4635 159
rect 4631 149 4635 153
rect 4631 143 4635 147
rect 4631 137 4635 141
rect 4631 131 4635 135
rect 4631 125 4635 129
rect 4631 119 4635 123
rect 4631 113 4635 117
rect 4631 107 4635 111
rect 4631 101 4635 105
rect 4631 95 4635 99
rect 4631 89 4635 93
rect 4631 83 4635 87
rect 4631 77 4635 81
rect 4631 71 4635 75
rect 4631 65 4635 69
rect 4631 59 4635 63
rect 4631 53 4635 57
rect 4631 47 4635 51
rect 4631 41 4635 45
rect 4631 35 4635 39
rect 4631 29 4635 33
rect 4631 23 4635 27
rect 4631 17 4635 21
rect 4631 11 4635 15
rect 4631 5 4635 9
<< polysilicon >>
rect 371 505 4629 506
rect 371 501 673 505
rect 677 501 679 505
rect 683 501 685 505
rect 689 501 691 505
rect 695 501 697 505
rect 701 501 703 505
rect 707 501 709 505
rect 713 501 969 505
rect 973 501 975 505
rect 979 501 981 505
rect 985 501 987 505
rect 991 501 993 505
rect 997 501 999 505
rect 1003 501 1005 505
rect 1009 501 1147 505
rect 1151 501 1153 505
rect 1157 501 1159 505
rect 1163 501 1165 505
rect 1169 501 1171 505
rect 1175 501 1177 505
rect 1181 501 1183 505
rect 1187 501 1443 505
rect 1447 501 1449 505
rect 1453 501 1455 505
rect 1459 501 1461 505
rect 1465 501 1467 505
rect 1471 501 1473 505
rect 1477 501 1479 505
rect 1483 501 1621 505
rect 1625 501 1627 505
rect 1631 501 1633 505
rect 1637 501 1639 505
rect 1643 501 1645 505
rect 1649 501 1651 505
rect 1655 501 1657 505
rect 1661 501 1917 505
rect 1921 501 1923 505
rect 1927 501 1929 505
rect 1933 501 1935 505
rect 1939 501 1941 505
rect 1945 501 1947 505
rect 1951 501 1953 505
rect 1957 501 2095 505
rect 2099 501 2101 505
rect 2105 501 2107 505
rect 2111 501 2113 505
rect 2117 501 2119 505
rect 2123 501 2125 505
rect 2129 501 2131 505
rect 2135 501 2391 505
rect 2395 501 2397 505
rect 2401 501 2403 505
rect 2407 501 2409 505
rect 2413 501 2415 505
rect 2419 501 2421 505
rect 2425 501 2427 505
rect 2431 501 2569 505
rect 2573 501 2575 505
rect 2579 501 2581 505
rect 2585 501 2587 505
rect 2591 501 2593 505
rect 2597 501 2599 505
rect 2603 501 2605 505
rect 2609 501 2865 505
rect 2869 501 2871 505
rect 2875 501 2877 505
rect 2881 501 2883 505
rect 2887 501 2889 505
rect 2893 501 2895 505
rect 2899 501 2901 505
rect 2905 501 3043 505
rect 3047 501 3049 505
rect 3053 501 3055 505
rect 3059 501 3061 505
rect 3065 501 3067 505
rect 3071 501 3073 505
rect 3077 501 3079 505
rect 3083 501 3339 505
rect 3343 501 3345 505
rect 3349 501 3351 505
rect 3355 501 3357 505
rect 3361 501 3363 505
rect 3367 501 3369 505
rect 3373 501 3375 505
rect 3379 501 3517 505
rect 3521 501 3523 505
rect 3527 501 3529 505
rect 3533 501 3535 505
rect 3539 501 3541 505
rect 3545 501 3547 505
rect 3551 501 3553 505
rect 3557 501 3813 505
rect 3817 501 3819 505
rect 3823 501 3825 505
rect 3829 501 3831 505
rect 3835 501 3837 505
rect 3841 501 3843 505
rect 3847 501 3849 505
rect 3853 501 3991 505
rect 3995 501 3997 505
rect 4001 501 4003 505
rect 4007 501 4009 505
rect 4013 501 4015 505
rect 4019 501 4021 505
rect 4025 501 4027 505
rect 4031 501 4287 505
rect 4291 501 4293 505
rect 4297 501 4299 505
rect 4303 501 4305 505
rect 4309 501 4311 505
rect 4315 501 4317 505
rect 4321 501 4323 505
rect 4327 501 4629 505
rect 371 376 4629 501
rect 371 372 495 376
rect 499 372 501 376
rect 505 372 507 376
rect 511 372 513 376
rect 517 372 519 376
rect 523 372 525 376
rect 529 372 531 376
rect 535 372 673 376
rect 677 372 679 376
rect 683 372 685 376
rect 689 372 691 376
rect 695 372 697 376
rect 701 372 703 376
rect 707 372 709 376
rect 713 372 969 376
rect 973 372 975 376
rect 979 372 981 376
rect 985 372 987 376
rect 991 372 993 376
rect 997 372 999 376
rect 1003 372 1005 376
rect 1009 372 1147 376
rect 1151 372 1153 376
rect 1157 372 1159 376
rect 1163 372 1165 376
rect 1169 372 1171 376
rect 1175 372 1177 376
rect 1181 372 1183 376
rect 1187 372 1443 376
rect 1447 372 1449 376
rect 1453 372 1455 376
rect 1459 372 1461 376
rect 1465 372 1467 376
rect 1471 372 1473 376
rect 1477 372 1479 376
rect 1483 372 1621 376
rect 1625 372 1627 376
rect 1631 372 1633 376
rect 1637 372 1639 376
rect 1643 372 1645 376
rect 1649 372 1651 376
rect 1655 372 1657 376
rect 1661 372 1917 376
rect 1921 372 1923 376
rect 1927 372 1929 376
rect 1933 372 1935 376
rect 1939 372 1941 376
rect 1945 372 1947 376
rect 1951 372 1953 376
rect 1957 372 2095 376
rect 2099 372 2101 376
rect 2105 372 2107 376
rect 2111 372 2113 376
rect 2117 372 2119 376
rect 2123 372 2125 376
rect 2129 372 2131 376
rect 2135 372 2391 376
rect 2395 372 2397 376
rect 2401 372 2403 376
rect 2407 372 2409 376
rect 2413 372 2415 376
rect 2419 372 2421 376
rect 2425 372 2427 376
rect 2431 372 2569 376
rect 2573 372 2575 376
rect 2579 372 2581 376
rect 2585 372 2587 376
rect 2591 372 2593 376
rect 2597 372 2599 376
rect 2603 372 2605 376
rect 2609 372 2865 376
rect 2869 372 2871 376
rect 2875 372 2877 376
rect 2881 372 2883 376
rect 2887 372 2889 376
rect 2893 372 2895 376
rect 2899 372 2901 376
rect 2905 372 3043 376
rect 3047 372 3049 376
rect 3053 372 3055 376
rect 3059 372 3061 376
rect 3065 372 3067 376
rect 3071 372 3073 376
rect 3077 372 3079 376
rect 3083 372 3339 376
rect 3343 372 3345 376
rect 3349 372 3351 376
rect 3355 372 3357 376
rect 3361 372 3363 376
rect 3367 372 3369 376
rect 3373 372 3375 376
rect 3379 372 3517 376
rect 3521 372 3523 376
rect 3527 372 3529 376
rect 3533 372 3535 376
rect 3539 372 3541 376
rect 3545 372 3547 376
rect 3551 372 3553 376
rect 3557 372 3813 376
rect 3817 372 3819 376
rect 3823 372 3825 376
rect 3829 372 3831 376
rect 3835 372 3837 376
rect 3841 372 3843 376
rect 3847 372 3849 376
rect 3853 372 3991 376
rect 3995 372 3997 376
rect 4001 372 4003 376
rect 4007 372 4009 376
rect 4013 372 4015 376
rect 4019 372 4021 376
rect 4025 372 4027 376
rect 4031 372 4287 376
rect 4291 372 4293 376
rect 4297 372 4299 376
rect 4303 372 4305 376
rect 4309 372 4311 376
rect 4315 372 4317 376
rect 4321 372 4323 376
rect 4327 372 4465 376
rect 4469 372 4471 376
rect 4475 372 4477 376
rect 4481 372 4483 376
rect 4487 372 4489 376
rect 4493 372 4495 376
rect 4499 372 4501 376
rect 4505 372 4629 376
rect 371 371 4629 372
rect 2 362 363 363
rect 2 358 3 362
rect 7 358 323 362
rect 327 358 329 362
rect 333 358 335 362
rect 339 358 341 362
rect 345 358 347 362
rect 351 358 353 362
rect 357 358 363 362
rect 2 357 363 358
rect 2 356 358 357
rect 2 352 3 356
rect 7 353 358 356
rect 362 353 363 357
rect 7 352 363 353
rect 2 351 363 352
rect 2 350 358 351
rect 2 346 3 350
rect 7 347 358 350
rect 362 347 363 351
rect 7 346 363 347
rect 2 345 363 346
rect 2 344 358 345
rect 2 340 3 344
rect 7 341 358 344
rect 362 341 363 345
rect 7 340 363 341
rect 2 339 363 340
rect 2 338 358 339
rect 2 334 3 338
rect 7 335 358 338
rect 362 335 363 339
rect 7 334 363 335
rect 2 333 363 334
rect 2 332 358 333
rect 2 328 3 332
rect 7 329 358 332
rect 362 329 363 333
rect 7 328 363 329
rect 2 327 363 328
rect 2 326 358 327
rect 2 322 3 326
rect 7 323 358 326
rect 362 323 363 327
rect 7 322 363 323
rect 2 320 363 322
rect 2 316 3 320
rect 7 316 363 320
rect 2 310 363 316
rect 310 7 363 310
rect 310 3 316 7
rect 320 3 322 7
rect 326 3 328 7
rect 332 3 334 7
rect 338 3 340 7
rect 344 3 346 7
rect 350 3 352 7
rect 356 3 358 7
rect 362 3 363 7
rect 310 2 363 3
rect 4637 362 4998 363
rect 4637 358 4643 362
rect 4647 358 4649 362
rect 4653 358 4655 362
rect 4659 358 4661 362
rect 4665 358 4667 362
rect 4671 358 4673 362
rect 4677 358 4993 362
rect 4997 358 4998 362
rect 4637 357 4998 358
rect 4637 353 4638 357
rect 4642 356 4998 357
rect 4642 353 4993 356
rect 4637 352 4993 353
rect 4997 352 4998 356
rect 4637 351 4998 352
rect 4637 347 4638 351
rect 4642 350 4998 351
rect 4642 347 4993 350
rect 4637 346 4993 347
rect 4997 346 4998 350
rect 4637 345 4998 346
rect 4637 341 4638 345
rect 4642 344 4998 345
rect 4642 341 4993 344
rect 4637 340 4993 341
rect 4997 340 4998 344
rect 4637 339 4998 340
rect 4637 335 4638 339
rect 4642 338 4998 339
rect 4642 335 4993 338
rect 4637 334 4993 335
rect 4997 334 4998 338
rect 4637 333 4998 334
rect 4637 329 4638 333
rect 4642 332 4998 333
rect 4642 329 4993 332
rect 4637 328 4993 329
rect 4997 328 4998 332
rect 4637 327 4998 328
rect 4637 323 4638 327
rect 4642 326 4998 327
rect 4642 323 4993 326
rect 4637 322 4993 323
rect 4997 322 4998 326
rect 4637 320 4998 322
rect 4637 316 4993 320
rect 4997 316 4998 320
rect 4637 310 4998 316
rect 4637 7 4690 310
rect 4637 3 4638 7
rect 4642 3 4644 7
rect 4648 3 4650 7
rect 4654 3 4656 7
rect 4660 3 4662 7
rect 4666 3 4668 7
rect 4672 3 4674 7
rect 4678 3 4680 7
rect 4684 3 4690 7
rect 4637 2 4690 3
<< polycontact >>
rect 673 501 677 505
rect 679 501 683 505
rect 685 501 689 505
rect 691 501 695 505
rect 697 501 701 505
rect 703 501 707 505
rect 709 501 713 505
rect 969 501 973 505
rect 975 501 979 505
rect 981 501 985 505
rect 987 501 991 505
rect 993 501 997 505
rect 999 501 1003 505
rect 1005 501 1009 505
rect 1147 501 1151 505
rect 1153 501 1157 505
rect 1159 501 1163 505
rect 1165 501 1169 505
rect 1171 501 1175 505
rect 1177 501 1181 505
rect 1183 501 1187 505
rect 1443 501 1447 505
rect 1449 501 1453 505
rect 1455 501 1459 505
rect 1461 501 1465 505
rect 1467 501 1471 505
rect 1473 501 1477 505
rect 1479 501 1483 505
rect 1621 501 1625 505
rect 1627 501 1631 505
rect 1633 501 1637 505
rect 1639 501 1643 505
rect 1645 501 1649 505
rect 1651 501 1655 505
rect 1657 501 1661 505
rect 1917 501 1921 505
rect 1923 501 1927 505
rect 1929 501 1933 505
rect 1935 501 1939 505
rect 1941 501 1945 505
rect 1947 501 1951 505
rect 1953 501 1957 505
rect 2095 501 2099 505
rect 2101 501 2105 505
rect 2107 501 2111 505
rect 2113 501 2117 505
rect 2119 501 2123 505
rect 2125 501 2129 505
rect 2131 501 2135 505
rect 2391 501 2395 505
rect 2397 501 2401 505
rect 2403 501 2407 505
rect 2409 501 2413 505
rect 2415 501 2419 505
rect 2421 501 2425 505
rect 2427 501 2431 505
rect 2569 501 2573 505
rect 2575 501 2579 505
rect 2581 501 2585 505
rect 2587 501 2591 505
rect 2593 501 2597 505
rect 2599 501 2603 505
rect 2605 501 2609 505
rect 2865 501 2869 505
rect 2871 501 2875 505
rect 2877 501 2881 505
rect 2883 501 2887 505
rect 2889 501 2893 505
rect 2895 501 2899 505
rect 2901 501 2905 505
rect 3043 501 3047 505
rect 3049 501 3053 505
rect 3055 501 3059 505
rect 3061 501 3065 505
rect 3067 501 3071 505
rect 3073 501 3077 505
rect 3079 501 3083 505
rect 3339 501 3343 505
rect 3345 501 3349 505
rect 3351 501 3355 505
rect 3357 501 3361 505
rect 3363 501 3367 505
rect 3369 501 3373 505
rect 3375 501 3379 505
rect 3517 501 3521 505
rect 3523 501 3527 505
rect 3529 501 3533 505
rect 3535 501 3539 505
rect 3541 501 3545 505
rect 3547 501 3551 505
rect 3553 501 3557 505
rect 3813 501 3817 505
rect 3819 501 3823 505
rect 3825 501 3829 505
rect 3831 501 3835 505
rect 3837 501 3841 505
rect 3843 501 3847 505
rect 3849 501 3853 505
rect 3991 501 3995 505
rect 3997 501 4001 505
rect 4003 501 4007 505
rect 4009 501 4013 505
rect 4015 501 4019 505
rect 4021 501 4025 505
rect 4027 501 4031 505
rect 4287 501 4291 505
rect 4293 501 4297 505
rect 4299 501 4303 505
rect 4305 501 4309 505
rect 4311 501 4315 505
rect 4317 501 4321 505
rect 4323 501 4327 505
rect 495 372 499 376
rect 501 372 505 376
rect 507 372 511 376
rect 513 372 517 376
rect 519 372 523 376
rect 525 372 529 376
rect 531 372 535 376
rect 673 372 677 376
rect 679 372 683 376
rect 685 372 689 376
rect 691 372 695 376
rect 697 372 701 376
rect 703 372 707 376
rect 709 372 713 376
rect 969 372 973 376
rect 975 372 979 376
rect 981 372 985 376
rect 987 372 991 376
rect 993 372 997 376
rect 999 372 1003 376
rect 1005 372 1009 376
rect 1147 372 1151 376
rect 1153 372 1157 376
rect 1159 372 1163 376
rect 1165 372 1169 376
rect 1171 372 1175 376
rect 1177 372 1181 376
rect 1183 372 1187 376
rect 1443 372 1447 376
rect 1449 372 1453 376
rect 1455 372 1459 376
rect 1461 372 1465 376
rect 1467 372 1471 376
rect 1473 372 1477 376
rect 1479 372 1483 376
rect 1621 372 1625 376
rect 1627 372 1631 376
rect 1633 372 1637 376
rect 1639 372 1643 376
rect 1645 372 1649 376
rect 1651 372 1655 376
rect 1657 372 1661 376
rect 1917 372 1921 376
rect 1923 372 1927 376
rect 1929 372 1933 376
rect 1935 372 1939 376
rect 1941 372 1945 376
rect 1947 372 1951 376
rect 1953 372 1957 376
rect 2095 372 2099 376
rect 2101 372 2105 376
rect 2107 372 2111 376
rect 2113 372 2117 376
rect 2119 372 2123 376
rect 2125 372 2129 376
rect 2131 372 2135 376
rect 2391 372 2395 376
rect 2397 372 2401 376
rect 2403 372 2407 376
rect 2409 372 2413 376
rect 2415 372 2419 376
rect 2421 372 2425 376
rect 2427 372 2431 376
rect 2569 372 2573 376
rect 2575 372 2579 376
rect 2581 372 2585 376
rect 2587 372 2591 376
rect 2593 372 2597 376
rect 2599 372 2603 376
rect 2605 372 2609 376
rect 2865 372 2869 376
rect 2871 372 2875 376
rect 2877 372 2881 376
rect 2883 372 2887 376
rect 2889 372 2893 376
rect 2895 372 2899 376
rect 2901 372 2905 376
rect 3043 372 3047 376
rect 3049 372 3053 376
rect 3055 372 3059 376
rect 3061 372 3065 376
rect 3067 372 3071 376
rect 3073 372 3077 376
rect 3079 372 3083 376
rect 3339 372 3343 376
rect 3345 372 3349 376
rect 3351 372 3355 376
rect 3357 372 3361 376
rect 3363 372 3367 376
rect 3369 372 3373 376
rect 3375 372 3379 376
rect 3517 372 3521 376
rect 3523 372 3527 376
rect 3529 372 3533 376
rect 3535 372 3539 376
rect 3541 372 3545 376
rect 3547 372 3551 376
rect 3553 372 3557 376
rect 3813 372 3817 376
rect 3819 372 3823 376
rect 3825 372 3829 376
rect 3831 372 3835 376
rect 3837 372 3841 376
rect 3843 372 3847 376
rect 3849 372 3853 376
rect 3991 372 3995 376
rect 3997 372 4001 376
rect 4003 372 4007 376
rect 4009 372 4013 376
rect 4015 372 4019 376
rect 4021 372 4025 376
rect 4027 372 4031 376
rect 4287 372 4291 376
rect 4293 372 4297 376
rect 4299 372 4303 376
rect 4305 372 4309 376
rect 4311 372 4315 376
rect 4317 372 4321 376
rect 4323 372 4327 376
rect 4465 372 4469 376
rect 4471 372 4475 376
rect 4477 372 4481 376
rect 4483 372 4487 376
rect 4489 372 4493 376
rect 4495 372 4499 376
rect 4501 372 4505 376
rect 3 358 7 362
rect 323 358 327 362
rect 329 358 333 362
rect 335 358 339 362
rect 341 358 345 362
rect 347 358 351 362
rect 353 358 357 362
rect 3 352 7 356
rect 358 353 362 357
rect 3 346 7 350
rect 358 347 362 351
rect 3 340 7 344
rect 358 341 362 345
rect 3 334 7 338
rect 358 335 362 339
rect 3 328 7 332
rect 358 329 362 333
rect 3 322 7 326
rect 358 323 362 327
rect 3 316 7 320
rect 316 3 320 7
rect 322 3 326 7
rect 328 3 332 7
rect 334 3 338 7
rect 340 3 344 7
rect 346 3 350 7
rect 352 3 356 7
rect 358 3 362 7
rect 4643 358 4647 362
rect 4649 358 4653 362
rect 4655 358 4659 362
rect 4661 358 4665 362
rect 4667 358 4671 362
rect 4673 358 4677 362
rect 4993 358 4997 362
rect 4638 353 4642 357
rect 4993 352 4997 356
rect 4638 347 4642 351
rect 4993 346 4997 350
rect 4638 341 4642 345
rect 4993 340 4997 344
rect 4638 335 4642 339
rect 4993 334 4997 338
rect 4638 329 4642 333
rect 4993 328 4997 332
rect 4638 323 4642 327
rect 4993 322 4997 326
rect 4993 316 4997 320
rect 4638 3 4642 7
rect 4644 3 4648 7
rect 4650 3 4654 7
rect 4656 3 4660 7
rect 4662 3 4666 7
rect 4668 3 4672 7
rect 4674 3 4678 7
rect 4680 3 4684 7
<< metal1 >>
rect 543 509 545 513
rect 549 509 551 513
rect 555 509 557 513
rect 561 509 563 513
rect 567 509 569 513
rect 573 509 575 513
rect 539 499 579 509
rect 543 495 545 499
rect 549 495 551 499
rect 555 495 557 499
rect 561 495 563 499
rect 567 495 569 499
rect 573 495 575 499
rect 539 493 579 495
rect 543 489 545 493
rect 549 489 551 493
rect 555 489 557 493
rect 561 489 563 493
rect 567 489 569 493
rect 573 489 575 493
rect 539 487 579 489
rect 543 483 545 487
rect 549 483 551 487
rect 555 483 557 487
rect 561 483 563 487
rect 567 483 569 487
rect 573 483 575 487
rect 539 481 579 483
rect 543 477 545 481
rect 549 477 551 481
rect 555 477 557 481
rect 561 477 563 481
rect 567 477 569 481
rect 573 477 575 481
rect 539 475 579 477
rect 543 471 545 475
rect 549 471 551 475
rect 555 471 557 475
rect 561 471 563 475
rect 567 471 569 475
rect 573 471 575 475
rect 539 470 579 471
rect 543 466 545 470
rect 549 466 551 470
rect 555 466 557 470
rect 561 466 563 470
rect 567 466 569 470
rect 573 466 575 470
rect 539 465 579 466
rect 495 450 535 451
rect 499 441 501 450
rect 505 441 507 450
rect 511 441 513 450
rect 517 441 519 450
rect 523 441 525 450
rect 529 441 531 450
rect 495 439 535 441
rect 499 435 501 439
rect 505 435 507 439
rect 511 435 513 439
rect 517 435 519 439
rect 523 435 525 439
rect 529 435 531 439
rect 495 433 535 435
rect 499 429 501 433
rect 505 429 507 433
rect 511 429 513 433
rect 517 429 519 433
rect 523 429 525 433
rect 529 429 531 433
rect 495 427 535 429
rect 499 423 501 427
rect 505 423 507 427
rect 511 423 513 427
rect 517 423 519 427
rect 523 423 525 427
rect 529 423 531 427
rect 495 421 535 423
rect 499 412 501 421
rect 505 412 507 421
rect 511 412 513 421
rect 517 412 519 421
rect 523 412 525 421
rect 529 412 531 421
rect 539 449 569 465
rect 583 461 592 509
rect 573 460 592 461
rect 577 456 578 460
rect 582 456 583 460
rect 587 456 588 460
rect 573 455 592 456
rect 616 461 625 509
rect 633 509 635 513
rect 639 509 641 513
rect 645 509 647 513
rect 651 509 653 513
rect 657 509 659 513
rect 663 509 665 513
rect 629 499 669 509
rect 633 495 635 499
rect 639 495 641 499
rect 645 495 647 499
rect 651 495 653 499
rect 657 495 659 499
rect 663 495 669 499
rect 629 493 669 495
rect 633 489 635 493
rect 639 489 641 493
rect 645 489 647 493
rect 651 489 653 493
rect 657 489 659 493
rect 663 489 665 493
rect 629 487 669 489
rect 633 483 635 487
rect 639 483 641 487
rect 645 483 647 487
rect 651 483 653 487
rect 657 483 659 487
rect 663 483 665 487
rect 629 481 669 483
rect 633 477 635 481
rect 639 477 641 481
rect 645 477 647 481
rect 651 477 653 481
rect 657 477 659 481
rect 663 477 665 481
rect 629 475 669 477
rect 633 471 635 475
rect 639 471 641 475
rect 645 471 647 475
rect 651 471 653 475
rect 657 471 659 475
rect 663 471 665 475
rect 629 470 669 471
rect 633 466 635 470
rect 639 466 641 470
rect 645 466 647 470
rect 651 466 653 470
rect 657 466 659 470
rect 663 466 665 470
rect 629 465 669 466
rect 616 460 635 461
rect 620 456 621 460
rect 625 456 626 460
rect 630 456 631 460
rect 616 455 635 456
rect 539 445 540 449
rect 544 445 546 449
rect 550 445 552 449
rect 556 445 558 449
rect 562 445 564 449
rect 568 445 569 449
rect 539 443 569 445
rect 539 439 540 443
rect 544 439 546 443
rect 550 439 552 443
rect 556 439 558 443
rect 562 439 564 443
rect 568 439 569 443
rect 539 437 569 439
rect 539 433 540 437
rect 544 433 546 437
rect 550 433 552 437
rect 556 433 558 437
rect 562 433 564 437
rect 568 433 569 437
rect 539 431 569 433
rect 539 427 540 431
rect 544 427 546 431
rect 550 427 552 431
rect 556 427 558 431
rect 562 427 564 431
rect 568 427 569 431
rect 539 424 569 427
rect 539 420 540 424
rect 544 420 546 424
rect 550 420 552 424
rect 556 420 558 424
rect 562 420 564 424
rect 568 420 569 424
rect 539 418 569 420
rect 539 414 540 418
rect 544 414 546 418
rect 550 414 552 418
rect 556 414 558 418
rect 562 414 564 418
rect 568 414 569 418
rect 539 413 569 414
rect 639 449 669 465
rect 639 445 640 449
rect 644 445 646 449
rect 650 445 652 449
rect 656 445 658 449
rect 662 445 664 449
rect 668 445 669 449
rect 639 443 669 445
rect 639 439 640 443
rect 644 439 646 443
rect 650 439 652 443
rect 656 439 658 443
rect 662 439 664 443
rect 668 439 669 443
rect 639 437 669 439
rect 639 433 640 437
rect 644 433 646 437
rect 650 433 652 437
rect 656 433 658 437
rect 662 433 664 437
rect 668 433 669 437
rect 639 431 669 433
rect 639 427 640 431
rect 644 427 646 431
rect 650 427 652 431
rect 656 427 658 431
rect 662 427 664 431
rect 668 427 669 431
rect 639 424 669 427
rect 639 420 640 424
rect 644 420 646 424
rect 650 420 652 424
rect 656 420 658 424
rect 662 420 664 424
rect 668 420 669 424
rect 639 418 669 420
rect 639 414 640 418
rect 644 414 646 418
rect 650 414 652 418
rect 656 414 658 418
rect 662 414 664 418
rect 668 414 669 418
rect 639 413 669 414
rect 677 509 679 513
rect 683 509 685 513
rect 689 509 691 513
rect 695 509 697 513
rect 701 509 703 513
rect 707 509 709 513
rect 673 505 713 509
rect 677 501 679 505
rect 683 501 685 505
rect 689 501 691 505
rect 695 501 697 505
rect 701 501 703 505
rect 707 501 709 505
rect 673 450 713 501
rect 677 441 679 450
rect 683 441 685 450
rect 689 441 691 450
rect 695 441 697 450
rect 701 441 703 450
rect 707 441 709 450
rect 673 439 713 441
rect 677 435 679 439
rect 683 435 685 439
rect 689 435 691 439
rect 695 435 697 439
rect 701 435 703 439
rect 707 435 709 439
rect 673 433 713 435
rect 677 429 679 433
rect 683 429 685 433
rect 689 429 691 433
rect 695 429 697 433
rect 701 429 703 433
rect 707 429 709 433
rect 673 427 713 429
rect 677 423 679 427
rect 683 423 685 427
rect 689 423 691 427
rect 695 423 697 427
rect 701 423 703 427
rect 707 423 709 427
rect 673 421 713 423
rect 495 376 535 412
rect 677 412 679 421
rect 683 412 685 421
rect 689 412 691 421
rect 695 412 697 421
rect 701 412 703 421
rect 707 412 709 421
rect 543 402 545 406
rect 549 402 551 406
rect 555 402 557 406
rect 561 402 563 406
rect 567 402 569 406
rect 573 402 575 406
rect 539 401 579 402
rect 543 397 545 401
rect 549 397 551 401
rect 555 397 557 401
rect 561 397 563 401
rect 567 397 569 401
rect 573 397 575 401
rect 539 394 579 397
rect 543 390 545 394
rect 549 390 551 394
rect 555 390 557 394
rect 561 390 563 394
rect 567 390 569 394
rect 573 390 575 394
rect 539 388 579 390
rect 543 384 545 388
rect 549 384 551 388
rect 555 384 557 388
rect 561 384 563 388
rect 567 384 569 388
rect 573 384 575 388
rect 545 382 579 384
rect 549 378 551 382
rect 555 378 557 382
rect 561 378 563 382
rect 567 378 569 382
rect 573 378 575 382
rect 633 402 635 406
rect 639 402 641 406
rect 645 402 647 406
rect 651 402 653 406
rect 657 402 659 406
rect 663 402 665 406
rect 629 401 669 402
rect 633 397 635 401
rect 639 397 641 401
rect 645 397 647 401
rect 651 397 653 401
rect 657 397 659 401
rect 663 397 665 401
rect 629 394 669 397
rect 633 390 635 394
rect 639 390 641 394
rect 645 390 647 394
rect 651 390 653 394
rect 657 390 659 394
rect 663 390 665 394
rect 629 388 669 390
rect 633 384 635 388
rect 639 384 641 388
rect 645 384 647 388
rect 651 384 653 388
rect 657 384 659 388
rect 663 384 665 388
rect 629 382 663 384
rect 633 378 635 382
rect 639 378 641 382
rect 645 378 647 382
rect 651 378 653 382
rect 657 378 659 382
rect 499 372 501 376
rect 505 372 507 376
rect 511 372 513 376
rect 517 372 519 376
rect 523 372 525 376
rect 529 372 531 376
rect 495 369 535 372
rect 673 376 713 412
rect 677 372 679 376
rect 683 372 685 376
rect 689 372 691 376
rect 695 372 697 376
rect 701 372 703 376
rect 707 372 709 376
rect 673 369 713 372
rect 973 509 975 513
rect 979 509 981 513
rect 985 509 987 513
rect 991 509 993 513
rect 997 509 999 513
rect 1003 509 1005 513
rect 969 505 1009 509
rect 973 501 975 505
rect 979 501 981 505
rect 985 501 987 505
rect 991 501 993 505
rect 997 501 999 505
rect 1003 501 1005 505
rect 969 450 1009 501
rect 973 441 975 450
rect 979 441 981 450
rect 985 441 987 450
rect 991 441 993 450
rect 997 441 999 450
rect 1003 441 1005 450
rect 969 439 1009 441
rect 973 435 975 439
rect 979 435 981 439
rect 985 435 987 439
rect 991 435 993 439
rect 997 435 999 439
rect 1003 435 1005 439
rect 969 433 1009 435
rect 973 429 975 433
rect 979 429 981 433
rect 985 429 987 433
rect 991 429 993 433
rect 997 429 999 433
rect 1003 429 1005 433
rect 969 427 1009 429
rect 973 423 975 427
rect 979 423 981 427
rect 985 423 987 427
rect 991 423 993 427
rect 997 423 999 427
rect 1003 423 1005 427
rect 969 421 1009 423
rect 973 412 975 421
rect 979 412 981 421
rect 985 412 987 421
rect 991 412 993 421
rect 997 412 999 421
rect 1003 412 1005 421
rect 1017 509 1019 513
rect 1023 509 1025 513
rect 1029 509 1031 513
rect 1035 509 1037 513
rect 1041 509 1043 513
rect 1047 509 1049 513
rect 1013 499 1053 509
rect 1013 495 1019 499
rect 1023 495 1025 499
rect 1029 495 1031 499
rect 1035 495 1037 499
rect 1041 495 1043 499
rect 1047 495 1049 499
rect 1013 493 1053 495
rect 1017 489 1019 493
rect 1023 489 1025 493
rect 1029 489 1031 493
rect 1035 489 1037 493
rect 1041 489 1043 493
rect 1047 489 1049 493
rect 1013 487 1053 489
rect 1017 483 1019 487
rect 1023 483 1025 487
rect 1029 483 1031 487
rect 1035 483 1037 487
rect 1041 483 1043 487
rect 1047 483 1049 487
rect 1013 481 1053 483
rect 1017 477 1019 481
rect 1023 477 1025 481
rect 1029 477 1031 481
rect 1035 477 1037 481
rect 1041 477 1043 481
rect 1047 477 1049 481
rect 1013 475 1053 477
rect 1017 471 1019 475
rect 1023 471 1025 475
rect 1029 471 1031 475
rect 1035 471 1037 475
rect 1041 471 1043 475
rect 1047 471 1049 475
rect 1013 469 1053 471
rect 1017 465 1019 469
rect 1023 465 1025 469
rect 1029 465 1031 469
rect 1035 465 1037 469
rect 1041 465 1043 469
rect 1047 465 1049 469
rect 1013 449 1043 465
rect 1057 461 1066 509
rect 1047 460 1066 461
rect 1051 456 1052 460
rect 1056 456 1057 460
rect 1061 456 1062 460
rect 1047 455 1066 456
rect 1090 461 1099 509
rect 1107 509 1109 513
rect 1113 509 1115 513
rect 1119 509 1121 513
rect 1125 509 1127 513
rect 1131 509 1133 513
rect 1137 509 1139 513
rect 1103 499 1143 509
rect 1107 495 1109 499
rect 1113 495 1115 499
rect 1119 495 1121 499
rect 1125 495 1127 499
rect 1131 495 1133 499
rect 1137 495 1143 499
rect 1103 493 1143 495
rect 1107 489 1109 493
rect 1113 489 1115 493
rect 1119 489 1121 493
rect 1125 489 1127 493
rect 1131 489 1133 493
rect 1137 489 1139 493
rect 1103 487 1143 489
rect 1107 483 1109 487
rect 1113 483 1115 487
rect 1119 483 1121 487
rect 1125 483 1127 487
rect 1131 483 1133 487
rect 1137 483 1139 487
rect 1103 481 1143 483
rect 1107 477 1109 481
rect 1113 477 1115 481
rect 1119 477 1121 481
rect 1125 477 1127 481
rect 1131 477 1133 481
rect 1137 477 1139 481
rect 1103 475 1143 477
rect 1107 471 1109 475
rect 1113 471 1115 475
rect 1119 471 1121 475
rect 1125 471 1127 475
rect 1131 471 1133 475
rect 1137 471 1139 475
rect 1103 469 1143 471
rect 1107 465 1109 469
rect 1113 465 1115 469
rect 1119 465 1121 469
rect 1125 465 1127 469
rect 1131 465 1133 469
rect 1137 465 1139 469
rect 1090 460 1109 461
rect 1094 456 1095 460
rect 1099 456 1100 460
rect 1104 456 1105 460
rect 1090 455 1109 456
rect 1013 445 1014 449
rect 1018 445 1020 449
rect 1024 445 1026 449
rect 1030 445 1032 449
rect 1036 445 1038 449
rect 1042 445 1043 449
rect 1013 443 1043 445
rect 1013 439 1014 443
rect 1018 439 1020 443
rect 1024 439 1026 443
rect 1030 439 1032 443
rect 1036 439 1038 443
rect 1042 439 1043 443
rect 1013 437 1043 439
rect 1013 433 1014 437
rect 1018 433 1020 437
rect 1024 433 1026 437
rect 1030 433 1032 437
rect 1036 433 1038 437
rect 1042 433 1043 437
rect 1013 431 1043 433
rect 1013 427 1014 431
rect 1018 427 1020 431
rect 1024 427 1026 431
rect 1030 427 1032 431
rect 1036 427 1038 431
rect 1042 427 1043 431
rect 1013 424 1043 427
rect 1013 420 1014 424
rect 1018 420 1020 424
rect 1024 420 1026 424
rect 1030 420 1032 424
rect 1036 420 1038 424
rect 1042 420 1043 424
rect 1013 418 1043 420
rect 1013 414 1014 418
rect 1018 414 1020 418
rect 1024 414 1026 418
rect 1030 414 1032 418
rect 1036 414 1038 418
rect 1042 414 1043 418
rect 1013 413 1043 414
rect 1113 449 1143 465
rect 1113 445 1114 449
rect 1118 445 1120 449
rect 1124 445 1126 449
rect 1130 445 1132 449
rect 1136 445 1138 449
rect 1142 445 1143 449
rect 1113 443 1143 445
rect 1113 439 1114 443
rect 1118 439 1120 443
rect 1124 439 1126 443
rect 1130 439 1132 443
rect 1136 439 1138 443
rect 1142 439 1143 443
rect 1113 437 1143 439
rect 1113 433 1114 437
rect 1118 433 1120 437
rect 1124 433 1126 437
rect 1130 433 1132 437
rect 1136 433 1138 437
rect 1142 433 1143 437
rect 1113 431 1143 433
rect 1113 427 1114 431
rect 1118 427 1120 431
rect 1124 427 1126 431
rect 1130 427 1132 431
rect 1136 427 1138 431
rect 1142 427 1143 431
rect 1113 424 1143 427
rect 1113 420 1114 424
rect 1118 420 1120 424
rect 1124 420 1126 424
rect 1130 420 1132 424
rect 1136 420 1138 424
rect 1142 420 1143 424
rect 1113 418 1143 420
rect 1113 414 1114 418
rect 1118 414 1120 418
rect 1124 414 1126 418
rect 1130 414 1132 418
rect 1136 414 1138 418
rect 1142 414 1143 418
rect 1113 413 1143 414
rect 1151 509 1153 513
rect 1157 509 1159 513
rect 1163 509 1165 513
rect 1169 509 1171 513
rect 1175 509 1177 513
rect 1181 509 1183 513
rect 1147 505 1187 509
rect 1151 501 1153 505
rect 1157 501 1159 505
rect 1163 501 1165 505
rect 1169 501 1171 505
rect 1175 501 1177 505
rect 1181 501 1183 505
rect 1147 450 1187 501
rect 1151 441 1153 450
rect 1157 441 1159 450
rect 1163 441 1165 450
rect 1169 441 1171 450
rect 1175 441 1177 450
rect 1181 441 1183 450
rect 1147 439 1187 441
rect 1151 435 1153 439
rect 1157 435 1159 439
rect 1163 435 1165 439
rect 1169 435 1171 439
rect 1175 435 1177 439
rect 1181 435 1183 439
rect 1147 433 1187 435
rect 1151 429 1153 433
rect 1157 429 1159 433
rect 1163 429 1165 433
rect 1169 429 1171 433
rect 1175 429 1177 433
rect 1181 429 1183 433
rect 1147 427 1187 429
rect 1151 423 1153 427
rect 1157 423 1159 427
rect 1163 423 1165 427
rect 1169 423 1171 427
rect 1175 423 1177 427
rect 1181 423 1183 427
rect 1147 421 1187 423
rect 969 376 1009 412
rect 1151 412 1153 421
rect 1157 412 1159 421
rect 1163 412 1165 421
rect 1169 412 1171 421
rect 1175 412 1177 421
rect 1181 412 1183 421
rect 1017 402 1019 406
rect 1023 402 1025 406
rect 1029 402 1031 406
rect 1035 402 1037 406
rect 1041 402 1043 406
rect 1047 402 1049 406
rect 1013 401 1053 402
rect 1017 397 1019 401
rect 1023 397 1025 401
rect 1029 397 1031 401
rect 1035 397 1037 401
rect 1041 397 1043 401
rect 1047 397 1049 401
rect 1013 394 1053 397
rect 1017 390 1019 394
rect 1023 390 1025 394
rect 1029 390 1031 394
rect 1035 390 1037 394
rect 1041 390 1043 394
rect 1047 390 1049 394
rect 1013 388 1053 390
rect 1017 384 1019 388
rect 1023 384 1025 388
rect 1029 384 1031 388
rect 1035 384 1037 388
rect 1041 384 1043 388
rect 1047 384 1049 388
rect 1019 382 1053 384
rect 1023 378 1025 382
rect 1029 378 1031 382
rect 1035 378 1037 382
rect 1041 378 1043 382
rect 1047 378 1049 382
rect 1107 402 1109 406
rect 1113 402 1115 406
rect 1119 402 1121 406
rect 1125 402 1127 406
rect 1131 402 1133 406
rect 1137 402 1139 406
rect 1103 401 1143 402
rect 1107 397 1109 401
rect 1113 397 1115 401
rect 1119 397 1121 401
rect 1125 397 1127 401
rect 1131 397 1133 401
rect 1137 397 1139 401
rect 1103 394 1143 397
rect 1107 390 1109 394
rect 1113 390 1115 394
rect 1119 390 1121 394
rect 1125 390 1127 394
rect 1131 390 1133 394
rect 1137 390 1139 394
rect 1103 388 1143 390
rect 1107 384 1109 388
rect 1113 384 1115 388
rect 1119 384 1121 388
rect 1125 384 1127 388
rect 1131 384 1133 388
rect 1137 384 1139 388
rect 1103 382 1137 384
rect 1107 378 1109 382
rect 1113 378 1115 382
rect 1119 378 1121 382
rect 1125 378 1127 382
rect 1131 378 1133 382
rect 973 372 975 376
rect 979 372 981 376
rect 985 372 987 376
rect 991 372 993 376
rect 997 372 999 376
rect 1003 372 1005 376
rect 969 369 1009 372
rect 1147 376 1187 412
rect 1151 372 1153 376
rect 1157 372 1159 376
rect 1163 372 1165 376
rect 1169 372 1171 376
rect 1175 372 1177 376
rect 1181 372 1183 376
rect 1147 369 1187 372
rect 1447 509 1449 513
rect 1453 509 1455 513
rect 1459 509 1461 513
rect 1465 509 1467 513
rect 1471 509 1473 513
rect 1477 509 1479 513
rect 1443 505 1483 509
rect 1447 501 1449 505
rect 1453 501 1455 505
rect 1459 501 1461 505
rect 1465 501 1467 505
rect 1471 501 1473 505
rect 1477 501 1479 505
rect 1443 450 1483 501
rect 1447 441 1449 450
rect 1453 441 1455 450
rect 1459 441 1461 450
rect 1465 441 1467 450
rect 1471 441 1473 450
rect 1477 441 1479 450
rect 1443 439 1483 441
rect 1447 435 1449 439
rect 1453 435 1455 439
rect 1459 435 1461 439
rect 1465 435 1467 439
rect 1471 435 1473 439
rect 1477 435 1479 439
rect 1443 433 1483 435
rect 1447 429 1449 433
rect 1453 429 1455 433
rect 1459 429 1461 433
rect 1465 429 1467 433
rect 1471 429 1473 433
rect 1477 429 1479 433
rect 1443 427 1483 429
rect 1447 423 1449 427
rect 1453 423 1455 427
rect 1459 423 1461 427
rect 1465 423 1467 427
rect 1471 423 1473 427
rect 1477 423 1479 427
rect 1443 421 1483 423
rect 1447 412 1449 421
rect 1453 412 1455 421
rect 1459 412 1461 421
rect 1465 412 1467 421
rect 1471 412 1473 421
rect 1477 412 1479 421
rect 1491 509 1493 513
rect 1497 509 1499 513
rect 1503 509 1505 513
rect 1509 509 1511 513
rect 1515 509 1517 513
rect 1521 509 1523 513
rect 1487 499 1527 509
rect 1487 495 1493 499
rect 1497 495 1499 499
rect 1503 495 1505 499
rect 1509 495 1511 499
rect 1515 495 1517 499
rect 1521 495 1523 499
rect 1487 493 1527 495
rect 1491 489 1493 493
rect 1497 489 1499 493
rect 1503 489 1505 493
rect 1509 489 1511 493
rect 1515 489 1517 493
rect 1521 489 1523 493
rect 1487 487 1527 489
rect 1491 483 1493 487
rect 1497 483 1499 487
rect 1503 483 1505 487
rect 1509 483 1511 487
rect 1515 483 1517 487
rect 1521 483 1523 487
rect 1487 481 1527 483
rect 1491 477 1493 481
rect 1497 477 1499 481
rect 1503 477 1505 481
rect 1509 477 1511 481
rect 1515 477 1517 481
rect 1521 477 1523 481
rect 1487 475 1527 477
rect 1491 471 1493 475
rect 1497 471 1499 475
rect 1503 471 1505 475
rect 1509 471 1511 475
rect 1515 471 1517 475
rect 1521 471 1523 475
rect 1487 469 1527 471
rect 1491 465 1493 469
rect 1497 465 1499 469
rect 1503 465 1505 469
rect 1509 465 1511 469
rect 1515 465 1517 469
rect 1521 465 1523 469
rect 1487 449 1517 465
rect 1531 461 1540 509
rect 1521 460 1540 461
rect 1525 456 1526 460
rect 1530 456 1531 460
rect 1535 456 1536 460
rect 1521 455 1540 456
rect 1564 461 1573 509
rect 1581 509 1583 513
rect 1587 509 1589 513
rect 1593 509 1595 513
rect 1599 509 1601 513
rect 1605 509 1607 513
rect 1611 509 1613 513
rect 1577 499 1617 509
rect 1581 495 1583 499
rect 1587 495 1589 499
rect 1593 495 1595 499
rect 1599 495 1601 499
rect 1605 495 1607 499
rect 1611 495 1617 499
rect 1577 493 1617 495
rect 1581 489 1583 493
rect 1587 489 1589 493
rect 1593 489 1595 493
rect 1599 489 1601 493
rect 1605 489 1607 493
rect 1611 489 1613 493
rect 1577 487 1617 489
rect 1581 483 1583 487
rect 1587 483 1589 487
rect 1593 483 1595 487
rect 1599 483 1601 487
rect 1605 483 1607 487
rect 1611 483 1613 487
rect 1577 481 1617 483
rect 1581 477 1583 481
rect 1587 477 1589 481
rect 1593 477 1595 481
rect 1599 477 1601 481
rect 1605 477 1607 481
rect 1611 477 1613 481
rect 1577 475 1617 477
rect 1581 471 1583 475
rect 1587 471 1589 475
rect 1593 471 1595 475
rect 1599 471 1601 475
rect 1605 471 1607 475
rect 1611 471 1613 475
rect 1577 469 1617 471
rect 1581 465 1583 469
rect 1587 465 1589 469
rect 1593 465 1595 469
rect 1599 465 1601 469
rect 1605 465 1607 469
rect 1611 465 1613 469
rect 1564 460 1583 461
rect 1568 456 1569 460
rect 1573 456 1574 460
rect 1578 456 1579 460
rect 1564 455 1583 456
rect 1487 445 1488 449
rect 1492 445 1494 449
rect 1498 445 1500 449
rect 1504 445 1506 449
rect 1510 445 1512 449
rect 1516 445 1517 449
rect 1487 443 1517 445
rect 1487 439 1488 443
rect 1492 439 1494 443
rect 1498 439 1500 443
rect 1504 439 1506 443
rect 1510 439 1512 443
rect 1516 439 1517 443
rect 1487 437 1517 439
rect 1487 433 1488 437
rect 1492 433 1494 437
rect 1498 433 1500 437
rect 1504 433 1506 437
rect 1510 433 1512 437
rect 1516 433 1517 437
rect 1487 431 1517 433
rect 1487 427 1488 431
rect 1492 427 1494 431
rect 1498 427 1500 431
rect 1504 427 1506 431
rect 1510 427 1512 431
rect 1516 427 1517 431
rect 1487 424 1517 427
rect 1487 420 1488 424
rect 1492 420 1494 424
rect 1498 420 1500 424
rect 1504 420 1506 424
rect 1510 420 1512 424
rect 1516 420 1517 424
rect 1487 418 1517 420
rect 1487 414 1488 418
rect 1492 414 1494 418
rect 1498 414 1500 418
rect 1504 414 1506 418
rect 1510 414 1512 418
rect 1516 414 1517 418
rect 1487 413 1517 414
rect 1587 449 1617 465
rect 1587 445 1588 449
rect 1592 445 1594 449
rect 1598 445 1600 449
rect 1604 445 1606 449
rect 1610 445 1612 449
rect 1616 445 1617 449
rect 1587 443 1617 445
rect 1587 439 1588 443
rect 1592 439 1594 443
rect 1598 439 1600 443
rect 1604 439 1606 443
rect 1610 439 1612 443
rect 1616 439 1617 443
rect 1587 437 1617 439
rect 1587 433 1588 437
rect 1592 433 1594 437
rect 1598 433 1600 437
rect 1604 433 1606 437
rect 1610 433 1612 437
rect 1616 433 1617 437
rect 1587 431 1617 433
rect 1587 427 1588 431
rect 1592 427 1594 431
rect 1598 427 1600 431
rect 1604 427 1606 431
rect 1610 427 1612 431
rect 1616 427 1617 431
rect 1587 424 1617 427
rect 1587 420 1588 424
rect 1592 420 1594 424
rect 1598 420 1600 424
rect 1604 420 1606 424
rect 1610 420 1612 424
rect 1616 420 1617 424
rect 1587 418 1617 420
rect 1587 414 1588 418
rect 1592 414 1594 418
rect 1598 414 1600 418
rect 1604 414 1606 418
rect 1610 414 1612 418
rect 1616 414 1617 418
rect 1587 413 1617 414
rect 1625 509 1627 513
rect 1631 509 1633 513
rect 1637 509 1639 513
rect 1643 509 1645 513
rect 1649 509 1651 513
rect 1655 509 1657 513
rect 1621 505 1661 509
rect 1625 501 1627 505
rect 1631 501 1633 505
rect 1637 501 1639 505
rect 1643 501 1645 505
rect 1649 501 1651 505
rect 1655 501 1657 505
rect 1621 450 1661 501
rect 1625 441 1627 450
rect 1631 441 1633 450
rect 1637 441 1639 450
rect 1643 441 1645 450
rect 1649 441 1651 450
rect 1655 441 1657 450
rect 1621 439 1661 441
rect 1625 435 1627 439
rect 1631 435 1633 439
rect 1637 435 1639 439
rect 1643 435 1645 439
rect 1649 435 1651 439
rect 1655 435 1657 439
rect 1621 433 1661 435
rect 1625 429 1627 433
rect 1631 429 1633 433
rect 1637 429 1639 433
rect 1643 429 1645 433
rect 1649 429 1651 433
rect 1655 429 1657 433
rect 1621 427 1661 429
rect 1625 423 1627 427
rect 1631 423 1633 427
rect 1637 423 1639 427
rect 1643 423 1645 427
rect 1649 423 1651 427
rect 1655 423 1657 427
rect 1621 421 1661 423
rect 1443 376 1483 412
rect 1625 412 1627 421
rect 1631 412 1633 421
rect 1637 412 1639 421
rect 1643 412 1645 421
rect 1649 412 1651 421
rect 1655 412 1657 421
rect 1491 402 1493 406
rect 1497 402 1499 406
rect 1503 402 1505 406
rect 1509 402 1511 406
rect 1515 402 1517 406
rect 1521 402 1523 406
rect 1487 401 1527 402
rect 1491 397 1493 401
rect 1497 397 1499 401
rect 1503 397 1505 401
rect 1509 397 1511 401
rect 1515 397 1517 401
rect 1521 397 1523 401
rect 1487 394 1527 397
rect 1491 390 1493 394
rect 1497 390 1499 394
rect 1503 390 1505 394
rect 1509 390 1511 394
rect 1515 390 1517 394
rect 1521 390 1523 394
rect 1487 388 1527 390
rect 1491 384 1493 388
rect 1497 384 1499 388
rect 1503 384 1505 388
rect 1509 384 1511 388
rect 1515 384 1517 388
rect 1521 384 1523 388
rect 1493 382 1527 384
rect 1497 378 1499 382
rect 1503 378 1505 382
rect 1509 378 1511 382
rect 1515 378 1517 382
rect 1521 378 1523 382
rect 1581 402 1583 406
rect 1587 402 1589 406
rect 1593 402 1595 406
rect 1599 402 1601 406
rect 1605 402 1607 406
rect 1611 402 1613 406
rect 1577 401 1617 402
rect 1581 397 1583 401
rect 1587 397 1589 401
rect 1593 397 1595 401
rect 1599 397 1601 401
rect 1605 397 1607 401
rect 1611 397 1613 401
rect 1577 394 1617 397
rect 1581 390 1583 394
rect 1587 390 1589 394
rect 1593 390 1595 394
rect 1599 390 1601 394
rect 1605 390 1607 394
rect 1611 390 1613 394
rect 1577 388 1617 390
rect 1581 384 1583 388
rect 1587 384 1589 388
rect 1593 384 1595 388
rect 1599 384 1601 388
rect 1605 384 1607 388
rect 1611 384 1613 388
rect 1577 382 1611 384
rect 1581 378 1583 382
rect 1587 378 1589 382
rect 1593 378 1595 382
rect 1599 378 1601 382
rect 1605 378 1607 382
rect 1447 372 1449 376
rect 1453 372 1455 376
rect 1459 372 1461 376
rect 1465 372 1467 376
rect 1471 372 1473 376
rect 1477 372 1479 376
rect 1443 369 1483 372
rect 1621 376 1661 412
rect 1625 372 1627 376
rect 1631 372 1633 376
rect 1637 372 1639 376
rect 1643 372 1645 376
rect 1649 372 1651 376
rect 1655 372 1657 376
rect 1621 369 1661 372
rect 1921 509 1923 513
rect 1927 509 1929 513
rect 1933 509 1935 513
rect 1939 509 1941 513
rect 1945 509 1947 513
rect 1951 509 1953 513
rect 1917 505 1957 509
rect 1921 501 1923 505
rect 1927 501 1929 505
rect 1933 501 1935 505
rect 1939 501 1941 505
rect 1945 501 1947 505
rect 1951 501 1953 505
rect 1917 450 1957 501
rect 1921 441 1923 450
rect 1927 441 1929 450
rect 1933 441 1935 450
rect 1939 441 1941 450
rect 1945 441 1947 450
rect 1951 441 1953 450
rect 1917 439 1957 441
rect 1921 435 1923 439
rect 1927 435 1929 439
rect 1933 435 1935 439
rect 1939 435 1941 439
rect 1945 435 1947 439
rect 1951 435 1953 439
rect 1917 433 1957 435
rect 1921 429 1923 433
rect 1927 429 1929 433
rect 1933 429 1935 433
rect 1939 429 1941 433
rect 1945 429 1947 433
rect 1951 429 1953 433
rect 1917 427 1957 429
rect 1921 423 1923 427
rect 1927 423 1929 427
rect 1933 423 1935 427
rect 1939 423 1941 427
rect 1945 423 1947 427
rect 1951 423 1953 427
rect 1917 421 1957 423
rect 1921 412 1923 421
rect 1927 412 1929 421
rect 1933 412 1935 421
rect 1939 412 1941 421
rect 1945 412 1947 421
rect 1951 412 1953 421
rect 1965 509 1967 513
rect 1971 509 1973 513
rect 1977 509 1979 513
rect 1983 509 1985 513
rect 1989 509 1991 513
rect 1995 509 1997 513
rect 1961 499 2001 509
rect 1961 495 1967 499
rect 1971 495 1973 499
rect 1977 495 1979 499
rect 1983 495 1985 499
rect 1989 495 1991 499
rect 1995 495 1997 499
rect 1961 493 2001 495
rect 1965 489 1967 493
rect 1971 489 1973 493
rect 1977 489 1979 493
rect 1983 489 1985 493
rect 1989 489 1991 493
rect 1995 489 1997 493
rect 1961 487 2001 489
rect 1965 483 1967 487
rect 1971 483 1973 487
rect 1977 483 1979 487
rect 1983 483 1985 487
rect 1989 483 1991 487
rect 1995 483 1997 487
rect 1961 481 2001 483
rect 1965 477 1967 481
rect 1971 477 1973 481
rect 1977 477 1979 481
rect 1983 477 1985 481
rect 1989 477 1991 481
rect 1995 477 1997 481
rect 1961 475 2001 477
rect 1965 471 1967 475
rect 1971 471 1973 475
rect 1977 471 1979 475
rect 1983 471 1985 475
rect 1989 471 1991 475
rect 1995 471 1997 475
rect 1961 469 2001 471
rect 1965 465 1967 469
rect 1971 465 1973 469
rect 1977 465 1979 469
rect 1983 465 1985 469
rect 1989 465 1991 469
rect 1995 465 1997 469
rect 1961 449 1991 465
rect 2005 461 2014 509
rect 1995 460 2014 461
rect 1999 456 2000 460
rect 2004 456 2005 460
rect 2009 456 2010 460
rect 1995 455 2014 456
rect 2038 461 2047 509
rect 2055 509 2057 513
rect 2061 509 2063 513
rect 2067 509 2069 513
rect 2073 509 2075 513
rect 2079 509 2081 513
rect 2085 509 2087 513
rect 2051 499 2091 509
rect 2055 495 2057 499
rect 2061 495 2063 499
rect 2067 495 2069 499
rect 2073 495 2075 499
rect 2079 495 2081 499
rect 2085 495 2091 499
rect 2051 493 2091 495
rect 2055 489 2057 493
rect 2061 489 2063 493
rect 2067 489 2069 493
rect 2073 489 2075 493
rect 2079 489 2081 493
rect 2085 489 2087 493
rect 2051 487 2091 489
rect 2055 483 2057 487
rect 2061 483 2063 487
rect 2067 483 2069 487
rect 2073 483 2075 487
rect 2079 483 2081 487
rect 2085 483 2087 487
rect 2051 481 2091 483
rect 2055 477 2057 481
rect 2061 477 2063 481
rect 2067 477 2069 481
rect 2073 477 2075 481
rect 2079 477 2081 481
rect 2085 477 2087 481
rect 2051 475 2091 477
rect 2055 471 2057 475
rect 2061 471 2063 475
rect 2067 471 2069 475
rect 2073 471 2075 475
rect 2079 471 2081 475
rect 2085 471 2087 475
rect 2051 469 2091 471
rect 2055 465 2057 469
rect 2061 465 2063 469
rect 2067 465 2069 469
rect 2073 465 2075 469
rect 2079 465 2081 469
rect 2085 465 2087 469
rect 2038 460 2057 461
rect 2042 456 2043 460
rect 2047 456 2048 460
rect 2052 456 2053 460
rect 2038 455 2057 456
rect 1961 445 1962 449
rect 1966 445 1968 449
rect 1972 445 1974 449
rect 1978 445 1980 449
rect 1984 445 1986 449
rect 1990 445 1991 449
rect 1961 443 1991 445
rect 1961 439 1962 443
rect 1966 439 1968 443
rect 1972 439 1974 443
rect 1978 439 1980 443
rect 1984 439 1986 443
rect 1990 439 1991 443
rect 1961 437 1991 439
rect 1961 433 1962 437
rect 1966 433 1968 437
rect 1972 433 1974 437
rect 1978 433 1980 437
rect 1984 433 1986 437
rect 1990 433 1991 437
rect 1961 431 1991 433
rect 1961 427 1962 431
rect 1966 427 1968 431
rect 1972 427 1974 431
rect 1978 427 1980 431
rect 1984 427 1986 431
rect 1990 427 1991 431
rect 1961 424 1991 427
rect 1961 420 1962 424
rect 1966 420 1968 424
rect 1972 420 1974 424
rect 1978 420 1980 424
rect 1984 420 1986 424
rect 1990 420 1991 424
rect 1961 418 1991 420
rect 1961 414 1962 418
rect 1966 414 1968 418
rect 1972 414 1974 418
rect 1978 414 1980 418
rect 1984 414 1986 418
rect 1990 414 1991 418
rect 1961 413 1991 414
rect 2061 449 2091 465
rect 2061 445 2062 449
rect 2066 445 2068 449
rect 2072 445 2074 449
rect 2078 445 2080 449
rect 2084 445 2086 449
rect 2090 445 2091 449
rect 2061 443 2091 445
rect 2061 439 2062 443
rect 2066 439 2068 443
rect 2072 439 2074 443
rect 2078 439 2080 443
rect 2084 439 2086 443
rect 2090 439 2091 443
rect 2061 437 2091 439
rect 2061 433 2062 437
rect 2066 433 2068 437
rect 2072 433 2074 437
rect 2078 433 2080 437
rect 2084 433 2086 437
rect 2090 433 2091 437
rect 2061 431 2091 433
rect 2061 427 2062 431
rect 2066 427 2068 431
rect 2072 427 2074 431
rect 2078 427 2080 431
rect 2084 427 2086 431
rect 2090 427 2091 431
rect 2061 424 2091 427
rect 2061 420 2062 424
rect 2066 420 2068 424
rect 2072 420 2074 424
rect 2078 420 2080 424
rect 2084 420 2086 424
rect 2090 420 2091 424
rect 2061 418 2091 420
rect 2061 414 2062 418
rect 2066 414 2068 418
rect 2072 414 2074 418
rect 2078 414 2080 418
rect 2084 414 2086 418
rect 2090 414 2091 418
rect 2061 413 2091 414
rect 2099 509 2101 513
rect 2105 509 2107 513
rect 2111 509 2113 513
rect 2117 509 2119 513
rect 2123 509 2125 513
rect 2129 509 2131 513
rect 2095 505 2135 509
rect 2099 501 2101 505
rect 2105 501 2107 505
rect 2111 501 2113 505
rect 2117 501 2119 505
rect 2123 501 2125 505
rect 2129 501 2131 505
rect 2095 450 2135 501
rect 2099 441 2101 450
rect 2105 441 2107 450
rect 2111 441 2113 450
rect 2117 441 2119 450
rect 2123 441 2125 450
rect 2129 441 2131 450
rect 2095 439 2135 441
rect 2099 435 2101 439
rect 2105 435 2107 439
rect 2111 435 2113 439
rect 2117 435 2119 439
rect 2123 435 2125 439
rect 2129 435 2131 439
rect 2095 433 2135 435
rect 2099 429 2101 433
rect 2105 429 2107 433
rect 2111 429 2113 433
rect 2117 429 2119 433
rect 2123 429 2125 433
rect 2129 429 2131 433
rect 2095 427 2135 429
rect 2099 423 2101 427
rect 2105 423 2107 427
rect 2111 423 2113 427
rect 2117 423 2119 427
rect 2123 423 2125 427
rect 2129 423 2131 427
rect 2095 421 2135 423
rect 1917 376 1957 412
rect 2099 412 2101 421
rect 2105 412 2107 421
rect 2111 412 2113 421
rect 2117 412 2119 421
rect 2123 412 2125 421
rect 2129 412 2131 421
rect 1965 402 1967 406
rect 1971 402 1973 406
rect 1977 402 1979 406
rect 1983 402 1985 406
rect 1989 402 1991 406
rect 1995 402 1997 406
rect 1961 401 2001 402
rect 1965 397 1967 401
rect 1971 397 1973 401
rect 1977 397 1979 401
rect 1983 397 1985 401
rect 1989 397 1991 401
rect 1995 397 1997 401
rect 1961 394 2001 397
rect 1965 390 1967 394
rect 1971 390 1973 394
rect 1977 390 1979 394
rect 1983 390 1985 394
rect 1989 390 1991 394
rect 1995 390 1997 394
rect 1961 388 2001 390
rect 1965 384 1967 388
rect 1971 384 1973 388
rect 1977 384 1979 388
rect 1983 384 1985 388
rect 1989 384 1991 388
rect 1995 384 1997 388
rect 1967 382 2001 384
rect 1971 378 1973 382
rect 1977 378 1979 382
rect 1983 378 1985 382
rect 1989 378 1991 382
rect 1995 378 1997 382
rect 2055 402 2057 406
rect 2061 402 2063 406
rect 2067 402 2069 406
rect 2073 402 2075 406
rect 2079 402 2081 406
rect 2085 402 2087 406
rect 2051 401 2091 402
rect 2055 397 2057 401
rect 2061 397 2063 401
rect 2067 397 2069 401
rect 2073 397 2075 401
rect 2079 397 2081 401
rect 2085 397 2087 401
rect 2051 394 2091 397
rect 2055 390 2057 394
rect 2061 390 2063 394
rect 2067 390 2069 394
rect 2073 390 2075 394
rect 2079 390 2081 394
rect 2085 390 2087 394
rect 2051 388 2091 390
rect 2055 384 2057 388
rect 2061 384 2063 388
rect 2067 384 2069 388
rect 2073 384 2075 388
rect 2079 384 2081 388
rect 2085 384 2087 388
rect 2051 382 2085 384
rect 2055 378 2057 382
rect 2061 378 2063 382
rect 2067 378 2069 382
rect 2073 378 2075 382
rect 2079 378 2081 382
rect 1921 372 1923 376
rect 1927 372 1929 376
rect 1933 372 1935 376
rect 1939 372 1941 376
rect 1945 372 1947 376
rect 1951 372 1953 376
rect 1917 369 1957 372
rect 2095 376 2135 412
rect 2099 372 2101 376
rect 2105 372 2107 376
rect 2111 372 2113 376
rect 2117 372 2119 376
rect 2123 372 2125 376
rect 2129 372 2131 376
rect 2095 369 2135 372
rect 2395 509 2397 513
rect 2401 509 2403 513
rect 2407 509 2409 513
rect 2413 509 2415 513
rect 2419 509 2421 513
rect 2425 509 2427 513
rect 2391 505 2431 509
rect 2395 501 2397 505
rect 2401 501 2403 505
rect 2407 501 2409 505
rect 2413 501 2415 505
rect 2419 501 2421 505
rect 2425 501 2427 505
rect 2391 450 2431 501
rect 2395 441 2397 450
rect 2401 441 2403 450
rect 2407 441 2409 450
rect 2413 441 2415 450
rect 2419 441 2421 450
rect 2425 441 2427 450
rect 2391 439 2431 441
rect 2395 435 2397 439
rect 2401 435 2403 439
rect 2407 435 2409 439
rect 2413 435 2415 439
rect 2419 435 2421 439
rect 2425 435 2427 439
rect 2391 433 2431 435
rect 2395 429 2397 433
rect 2401 429 2403 433
rect 2407 429 2409 433
rect 2413 429 2415 433
rect 2419 429 2421 433
rect 2425 429 2427 433
rect 2391 427 2431 429
rect 2395 423 2397 427
rect 2401 423 2403 427
rect 2407 423 2409 427
rect 2413 423 2415 427
rect 2419 423 2421 427
rect 2425 423 2427 427
rect 2391 421 2431 423
rect 2395 412 2397 421
rect 2401 412 2403 421
rect 2407 412 2409 421
rect 2413 412 2415 421
rect 2419 412 2421 421
rect 2425 412 2427 421
rect 2439 509 2441 513
rect 2445 509 2447 513
rect 2451 509 2453 513
rect 2457 509 2459 513
rect 2463 509 2465 513
rect 2469 509 2471 513
rect 2435 499 2475 509
rect 2435 495 2441 499
rect 2445 495 2447 499
rect 2451 495 2453 499
rect 2457 495 2459 499
rect 2463 495 2465 499
rect 2469 495 2471 499
rect 2435 493 2475 495
rect 2439 489 2441 493
rect 2445 489 2447 493
rect 2451 489 2453 493
rect 2457 489 2459 493
rect 2463 489 2465 493
rect 2469 489 2471 493
rect 2435 487 2475 489
rect 2439 483 2441 487
rect 2445 483 2447 487
rect 2451 483 2453 487
rect 2457 483 2459 487
rect 2463 483 2465 487
rect 2469 483 2471 487
rect 2435 481 2475 483
rect 2439 477 2441 481
rect 2445 477 2447 481
rect 2451 477 2453 481
rect 2457 477 2459 481
rect 2463 477 2465 481
rect 2469 477 2471 481
rect 2435 475 2475 477
rect 2439 471 2441 475
rect 2445 471 2447 475
rect 2451 471 2453 475
rect 2457 471 2459 475
rect 2463 471 2465 475
rect 2469 471 2471 475
rect 2435 469 2475 471
rect 2439 465 2441 469
rect 2445 465 2447 469
rect 2451 465 2453 469
rect 2457 465 2459 469
rect 2463 465 2465 469
rect 2469 465 2471 469
rect 2435 449 2465 465
rect 2479 461 2488 509
rect 2469 460 2488 461
rect 2473 456 2474 460
rect 2478 456 2479 460
rect 2483 456 2484 460
rect 2469 455 2488 456
rect 2512 461 2521 509
rect 2529 509 2531 513
rect 2535 509 2537 513
rect 2541 509 2543 513
rect 2547 509 2549 513
rect 2553 509 2555 513
rect 2559 509 2561 513
rect 2525 499 2565 509
rect 2529 495 2531 499
rect 2535 495 2537 499
rect 2541 495 2543 499
rect 2547 495 2549 499
rect 2553 495 2555 499
rect 2559 495 2565 499
rect 2525 493 2565 495
rect 2529 489 2531 493
rect 2535 489 2537 493
rect 2541 489 2543 493
rect 2547 489 2549 493
rect 2553 489 2555 493
rect 2559 489 2561 493
rect 2525 487 2565 489
rect 2529 483 2531 487
rect 2535 483 2537 487
rect 2541 483 2543 487
rect 2547 483 2549 487
rect 2553 483 2555 487
rect 2559 483 2561 487
rect 2525 481 2565 483
rect 2529 477 2531 481
rect 2535 477 2537 481
rect 2541 477 2543 481
rect 2547 477 2549 481
rect 2553 477 2555 481
rect 2559 477 2561 481
rect 2525 475 2565 477
rect 2529 471 2531 475
rect 2535 471 2537 475
rect 2541 471 2543 475
rect 2547 471 2549 475
rect 2553 471 2555 475
rect 2559 471 2561 475
rect 2525 469 2565 471
rect 2529 465 2531 469
rect 2535 465 2537 469
rect 2541 465 2543 469
rect 2547 465 2549 469
rect 2553 465 2555 469
rect 2559 465 2561 469
rect 2512 460 2531 461
rect 2516 456 2517 460
rect 2521 456 2522 460
rect 2526 456 2527 460
rect 2512 455 2531 456
rect 2435 445 2436 449
rect 2440 445 2442 449
rect 2446 445 2448 449
rect 2452 445 2454 449
rect 2458 445 2460 449
rect 2464 445 2465 449
rect 2435 443 2465 445
rect 2435 439 2436 443
rect 2440 439 2442 443
rect 2446 439 2448 443
rect 2452 439 2454 443
rect 2458 439 2460 443
rect 2464 439 2465 443
rect 2435 437 2465 439
rect 2435 433 2436 437
rect 2440 433 2442 437
rect 2446 433 2448 437
rect 2452 433 2454 437
rect 2458 433 2460 437
rect 2464 433 2465 437
rect 2435 431 2465 433
rect 2435 427 2436 431
rect 2440 427 2442 431
rect 2446 427 2448 431
rect 2452 427 2454 431
rect 2458 427 2460 431
rect 2464 427 2465 431
rect 2435 424 2465 427
rect 2435 420 2436 424
rect 2440 420 2442 424
rect 2446 420 2448 424
rect 2452 420 2454 424
rect 2458 420 2460 424
rect 2464 420 2465 424
rect 2435 418 2465 420
rect 2435 414 2436 418
rect 2440 414 2442 418
rect 2446 414 2448 418
rect 2452 414 2454 418
rect 2458 414 2460 418
rect 2464 414 2465 418
rect 2435 413 2465 414
rect 2535 449 2565 465
rect 2535 445 2536 449
rect 2540 445 2542 449
rect 2546 445 2548 449
rect 2552 445 2554 449
rect 2558 445 2560 449
rect 2564 445 2565 449
rect 2535 443 2565 445
rect 2535 439 2536 443
rect 2540 439 2542 443
rect 2546 439 2548 443
rect 2552 439 2554 443
rect 2558 439 2560 443
rect 2564 439 2565 443
rect 2535 437 2565 439
rect 2535 433 2536 437
rect 2540 433 2542 437
rect 2546 433 2548 437
rect 2552 433 2554 437
rect 2558 433 2560 437
rect 2564 433 2565 437
rect 2535 431 2565 433
rect 2535 427 2536 431
rect 2540 427 2542 431
rect 2546 427 2548 431
rect 2552 427 2554 431
rect 2558 427 2560 431
rect 2564 427 2565 431
rect 2535 424 2565 427
rect 2535 420 2536 424
rect 2540 420 2542 424
rect 2546 420 2548 424
rect 2552 420 2554 424
rect 2558 420 2560 424
rect 2564 420 2565 424
rect 2535 418 2565 420
rect 2535 414 2536 418
rect 2540 414 2542 418
rect 2546 414 2548 418
rect 2552 414 2554 418
rect 2558 414 2560 418
rect 2564 414 2565 418
rect 2535 413 2565 414
rect 2573 509 2575 513
rect 2579 509 2581 513
rect 2585 509 2587 513
rect 2591 509 2593 513
rect 2597 509 2599 513
rect 2603 509 2605 513
rect 2569 505 2609 509
rect 2573 501 2575 505
rect 2579 501 2581 505
rect 2585 501 2587 505
rect 2591 501 2593 505
rect 2597 501 2599 505
rect 2603 501 2605 505
rect 2569 450 2609 501
rect 2573 441 2575 450
rect 2579 441 2581 450
rect 2585 441 2587 450
rect 2591 441 2593 450
rect 2597 441 2599 450
rect 2603 441 2605 450
rect 2569 439 2609 441
rect 2573 435 2575 439
rect 2579 435 2581 439
rect 2585 435 2587 439
rect 2591 435 2593 439
rect 2597 435 2599 439
rect 2603 435 2605 439
rect 2569 433 2609 435
rect 2573 429 2575 433
rect 2579 429 2581 433
rect 2585 429 2587 433
rect 2591 429 2593 433
rect 2597 429 2599 433
rect 2603 429 2605 433
rect 2569 427 2609 429
rect 2573 423 2575 427
rect 2579 423 2581 427
rect 2585 423 2587 427
rect 2591 423 2593 427
rect 2597 423 2599 427
rect 2603 423 2605 427
rect 2569 421 2609 423
rect 2391 376 2431 412
rect 2573 412 2575 421
rect 2579 412 2581 421
rect 2585 412 2587 421
rect 2591 412 2593 421
rect 2597 412 2599 421
rect 2603 412 2605 421
rect 2439 402 2441 406
rect 2445 402 2447 406
rect 2451 402 2453 406
rect 2457 402 2459 406
rect 2463 402 2465 406
rect 2469 402 2471 406
rect 2435 401 2475 402
rect 2439 397 2441 401
rect 2445 397 2447 401
rect 2451 397 2453 401
rect 2457 397 2459 401
rect 2463 397 2465 401
rect 2469 397 2471 401
rect 2435 394 2475 397
rect 2439 390 2441 394
rect 2445 390 2447 394
rect 2451 390 2453 394
rect 2457 390 2459 394
rect 2463 390 2465 394
rect 2469 390 2471 394
rect 2435 388 2475 390
rect 2439 384 2441 388
rect 2445 384 2447 388
rect 2451 384 2453 388
rect 2457 384 2459 388
rect 2463 384 2465 388
rect 2469 384 2471 388
rect 2441 382 2475 384
rect 2445 378 2447 382
rect 2451 378 2453 382
rect 2457 378 2459 382
rect 2463 378 2465 382
rect 2469 378 2471 382
rect 2529 402 2531 406
rect 2535 402 2537 406
rect 2541 402 2543 406
rect 2547 402 2549 406
rect 2553 402 2555 406
rect 2559 402 2561 406
rect 2525 401 2565 402
rect 2529 397 2531 401
rect 2535 397 2537 401
rect 2541 397 2543 401
rect 2547 397 2549 401
rect 2553 397 2555 401
rect 2559 397 2561 401
rect 2525 394 2565 397
rect 2529 390 2531 394
rect 2535 390 2537 394
rect 2541 390 2543 394
rect 2547 390 2549 394
rect 2553 390 2555 394
rect 2559 390 2561 394
rect 2525 388 2565 390
rect 2529 384 2531 388
rect 2535 384 2537 388
rect 2541 384 2543 388
rect 2547 384 2549 388
rect 2553 384 2555 388
rect 2559 384 2561 388
rect 2525 382 2559 384
rect 2529 378 2531 382
rect 2535 378 2537 382
rect 2541 378 2543 382
rect 2547 378 2549 382
rect 2553 378 2555 382
rect 2395 372 2397 376
rect 2401 372 2403 376
rect 2407 372 2409 376
rect 2413 372 2415 376
rect 2419 372 2421 376
rect 2425 372 2427 376
rect 2391 369 2431 372
rect 2569 376 2609 412
rect 2573 372 2575 376
rect 2579 372 2581 376
rect 2585 372 2587 376
rect 2591 372 2593 376
rect 2597 372 2599 376
rect 2603 372 2605 376
rect 2569 369 2609 372
rect 2869 509 2871 513
rect 2875 509 2877 513
rect 2881 509 2883 513
rect 2887 509 2889 513
rect 2893 509 2895 513
rect 2899 509 2901 513
rect 2865 505 2905 509
rect 2869 501 2871 505
rect 2875 501 2877 505
rect 2881 501 2883 505
rect 2887 501 2889 505
rect 2893 501 2895 505
rect 2899 501 2901 505
rect 2865 450 2905 501
rect 2869 441 2871 450
rect 2875 441 2877 450
rect 2881 441 2883 450
rect 2887 441 2889 450
rect 2893 441 2895 450
rect 2899 441 2901 450
rect 2865 439 2905 441
rect 2869 435 2871 439
rect 2875 435 2877 439
rect 2881 435 2883 439
rect 2887 435 2889 439
rect 2893 435 2895 439
rect 2899 435 2901 439
rect 2865 433 2905 435
rect 2869 429 2871 433
rect 2875 429 2877 433
rect 2881 429 2883 433
rect 2887 429 2889 433
rect 2893 429 2895 433
rect 2899 429 2901 433
rect 2865 427 2905 429
rect 2869 423 2871 427
rect 2875 423 2877 427
rect 2881 423 2883 427
rect 2887 423 2889 427
rect 2893 423 2895 427
rect 2899 423 2901 427
rect 2865 421 2905 423
rect 2869 412 2871 421
rect 2875 412 2877 421
rect 2881 412 2883 421
rect 2887 412 2889 421
rect 2893 412 2895 421
rect 2899 412 2901 421
rect 2913 509 2915 513
rect 2919 509 2921 513
rect 2925 509 2927 513
rect 2931 509 2933 513
rect 2937 509 2939 513
rect 2943 509 2945 513
rect 2909 499 2949 509
rect 2909 495 2915 499
rect 2919 495 2921 499
rect 2925 495 2927 499
rect 2931 495 2933 499
rect 2937 495 2939 499
rect 2943 495 2945 499
rect 2909 493 2949 495
rect 2913 489 2915 493
rect 2919 489 2921 493
rect 2925 489 2927 493
rect 2931 489 2933 493
rect 2937 489 2939 493
rect 2943 489 2945 493
rect 2909 487 2949 489
rect 2913 483 2915 487
rect 2919 483 2921 487
rect 2925 483 2927 487
rect 2931 483 2933 487
rect 2937 483 2939 487
rect 2943 483 2945 487
rect 2909 481 2949 483
rect 2913 477 2915 481
rect 2919 477 2921 481
rect 2925 477 2927 481
rect 2931 477 2933 481
rect 2937 477 2939 481
rect 2943 477 2945 481
rect 2909 475 2949 477
rect 2913 471 2915 475
rect 2919 471 2921 475
rect 2925 471 2927 475
rect 2931 471 2933 475
rect 2937 471 2939 475
rect 2943 471 2945 475
rect 2909 469 2949 471
rect 2913 465 2915 469
rect 2919 465 2921 469
rect 2925 465 2927 469
rect 2931 465 2933 469
rect 2937 465 2939 469
rect 2943 465 2945 469
rect 2909 449 2939 465
rect 2953 461 2962 509
rect 2943 460 2962 461
rect 2947 456 2948 460
rect 2952 456 2953 460
rect 2957 456 2958 460
rect 2943 455 2962 456
rect 2986 461 2995 509
rect 3003 509 3005 513
rect 3009 509 3011 513
rect 3015 509 3017 513
rect 3021 509 3023 513
rect 3027 509 3029 513
rect 3033 509 3035 513
rect 2999 499 3039 509
rect 3003 495 3005 499
rect 3009 495 3011 499
rect 3015 495 3017 499
rect 3021 495 3023 499
rect 3027 495 3029 499
rect 3033 495 3039 499
rect 2999 493 3039 495
rect 3003 489 3005 493
rect 3009 489 3011 493
rect 3015 489 3017 493
rect 3021 489 3023 493
rect 3027 489 3029 493
rect 3033 489 3035 493
rect 2999 487 3039 489
rect 3003 483 3005 487
rect 3009 483 3011 487
rect 3015 483 3017 487
rect 3021 483 3023 487
rect 3027 483 3029 487
rect 3033 483 3035 487
rect 2999 481 3039 483
rect 3003 477 3005 481
rect 3009 477 3011 481
rect 3015 477 3017 481
rect 3021 477 3023 481
rect 3027 477 3029 481
rect 3033 477 3035 481
rect 2999 475 3039 477
rect 3003 471 3005 475
rect 3009 471 3011 475
rect 3015 471 3017 475
rect 3021 471 3023 475
rect 3027 471 3029 475
rect 3033 471 3035 475
rect 2999 469 3039 471
rect 3003 465 3005 469
rect 3009 465 3011 469
rect 3015 465 3017 469
rect 3021 465 3023 469
rect 3027 465 3029 469
rect 3033 465 3035 469
rect 2986 460 3005 461
rect 2990 456 2991 460
rect 2995 456 2996 460
rect 3000 456 3001 460
rect 2986 455 3005 456
rect 2909 445 2910 449
rect 2914 445 2916 449
rect 2920 445 2922 449
rect 2926 445 2928 449
rect 2932 445 2934 449
rect 2938 445 2939 449
rect 2909 443 2939 445
rect 2909 439 2910 443
rect 2914 439 2916 443
rect 2920 439 2922 443
rect 2926 439 2928 443
rect 2932 439 2934 443
rect 2938 439 2939 443
rect 2909 437 2939 439
rect 2909 433 2910 437
rect 2914 433 2916 437
rect 2920 433 2922 437
rect 2926 433 2928 437
rect 2932 433 2934 437
rect 2938 433 2939 437
rect 2909 431 2939 433
rect 2909 427 2910 431
rect 2914 427 2916 431
rect 2920 427 2922 431
rect 2926 427 2928 431
rect 2932 427 2934 431
rect 2938 427 2939 431
rect 2909 424 2939 427
rect 2909 420 2910 424
rect 2914 420 2916 424
rect 2920 420 2922 424
rect 2926 420 2928 424
rect 2932 420 2934 424
rect 2938 420 2939 424
rect 2909 418 2939 420
rect 2909 414 2910 418
rect 2914 414 2916 418
rect 2920 414 2922 418
rect 2926 414 2928 418
rect 2932 414 2934 418
rect 2938 414 2939 418
rect 2909 413 2939 414
rect 3009 449 3039 465
rect 3009 445 3010 449
rect 3014 445 3016 449
rect 3020 445 3022 449
rect 3026 445 3028 449
rect 3032 445 3034 449
rect 3038 445 3039 449
rect 3009 443 3039 445
rect 3009 439 3010 443
rect 3014 439 3016 443
rect 3020 439 3022 443
rect 3026 439 3028 443
rect 3032 439 3034 443
rect 3038 439 3039 443
rect 3009 437 3039 439
rect 3009 433 3010 437
rect 3014 433 3016 437
rect 3020 433 3022 437
rect 3026 433 3028 437
rect 3032 433 3034 437
rect 3038 433 3039 437
rect 3009 431 3039 433
rect 3009 427 3010 431
rect 3014 427 3016 431
rect 3020 427 3022 431
rect 3026 427 3028 431
rect 3032 427 3034 431
rect 3038 427 3039 431
rect 3009 424 3039 427
rect 3009 420 3010 424
rect 3014 420 3016 424
rect 3020 420 3022 424
rect 3026 420 3028 424
rect 3032 420 3034 424
rect 3038 420 3039 424
rect 3009 418 3039 420
rect 3009 414 3010 418
rect 3014 414 3016 418
rect 3020 414 3022 418
rect 3026 414 3028 418
rect 3032 414 3034 418
rect 3038 414 3039 418
rect 3009 413 3039 414
rect 3047 509 3049 513
rect 3053 509 3055 513
rect 3059 509 3061 513
rect 3065 509 3067 513
rect 3071 509 3073 513
rect 3077 509 3079 513
rect 3043 505 3083 509
rect 3047 501 3049 505
rect 3053 501 3055 505
rect 3059 501 3061 505
rect 3065 501 3067 505
rect 3071 501 3073 505
rect 3077 501 3079 505
rect 3043 450 3083 501
rect 3047 441 3049 450
rect 3053 441 3055 450
rect 3059 441 3061 450
rect 3065 441 3067 450
rect 3071 441 3073 450
rect 3077 441 3079 450
rect 3043 439 3083 441
rect 3047 435 3049 439
rect 3053 435 3055 439
rect 3059 435 3061 439
rect 3065 435 3067 439
rect 3071 435 3073 439
rect 3077 435 3079 439
rect 3043 433 3083 435
rect 3047 429 3049 433
rect 3053 429 3055 433
rect 3059 429 3061 433
rect 3065 429 3067 433
rect 3071 429 3073 433
rect 3077 429 3079 433
rect 3043 427 3083 429
rect 3047 423 3049 427
rect 3053 423 3055 427
rect 3059 423 3061 427
rect 3065 423 3067 427
rect 3071 423 3073 427
rect 3077 423 3079 427
rect 3043 421 3083 423
rect 2865 376 2905 412
rect 3047 412 3049 421
rect 3053 412 3055 421
rect 3059 412 3061 421
rect 3065 412 3067 421
rect 3071 412 3073 421
rect 3077 412 3079 421
rect 2913 402 2915 406
rect 2919 402 2921 406
rect 2925 402 2927 406
rect 2931 402 2933 406
rect 2937 402 2939 406
rect 2943 402 2945 406
rect 2909 401 2949 402
rect 2913 397 2915 401
rect 2919 397 2921 401
rect 2925 397 2927 401
rect 2931 397 2933 401
rect 2937 397 2939 401
rect 2943 397 2945 401
rect 2909 394 2949 397
rect 2913 390 2915 394
rect 2919 390 2921 394
rect 2925 390 2927 394
rect 2931 390 2933 394
rect 2937 390 2939 394
rect 2943 390 2945 394
rect 2909 388 2949 390
rect 2913 384 2915 388
rect 2919 384 2921 388
rect 2925 384 2927 388
rect 2931 384 2933 388
rect 2937 384 2939 388
rect 2943 384 2945 388
rect 2915 382 2949 384
rect 2919 378 2921 382
rect 2925 378 2927 382
rect 2931 378 2933 382
rect 2937 378 2939 382
rect 2943 378 2945 382
rect 3003 402 3005 406
rect 3009 402 3011 406
rect 3015 402 3017 406
rect 3021 402 3023 406
rect 3027 402 3029 406
rect 3033 402 3035 406
rect 2999 401 3039 402
rect 3003 397 3005 401
rect 3009 397 3011 401
rect 3015 397 3017 401
rect 3021 397 3023 401
rect 3027 397 3029 401
rect 3033 397 3035 401
rect 2999 394 3039 397
rect 3003 390 3005 394
rect 3009 390 3011 394
rect 3015 390 3017 394
rect 3021 390 3023 394
rect 3027 390 3029 394
rect 3033 390 3035 394
rect 2999 388 3039 390
rect 3003 384 3005 388
rect 3009 384 3011 388
rect 3015 384 3017 388
rect 3021 384 3023 388
rect 3027 384 3029 388
rect 3033 384 3035 388
rect 2999 382 3033 384
rect 3003 378 3005 382
rect 3009 378 3011 382
rect 3015 378 3017 382
rect 3021 378 3023 382
rect 3027 378 3029 382
rect 2869 372 2871 376
rect 2875 372 2877 376
rect 2881 372 2883 376
rect 2887 372 2889 376
rect 2893 372 2895 376
rect 2899 372 2901 376
rect 2865 369 2905 372
rect 3043 376 3083 412
rect 3047 372 3049 376
rect 3053 372 3055 376
rect 3059 372 3061 376
rect 3065 372 3067 376
rect 3071 372 3073 376
rect 3077 372 3079 376
rect 3043 369 3083 372
rect 3343 509 3345 513
rect 3349 509 3351 513
rect 3355 509 3357 513
rect 3361 509 3363 513
rect 3367 509 3369 513
rect 3373 509 3375 513
rect 3339 505 3379 509
rect 3343 501 3345 505
rect 3349 501 3351 505
rect 3355 501 3357 505
rect 3361 501 3363 505
rect 3367 501 3369 505
rect 3373 501 3375 505
rect 3339 450 3379 501
rect 3343 441 3345 450
rect 3349 441 3351 450
rect 3355 441 3357 450
rect 3361 441 3363 450
rect 3367 441 3369 450
rect 3373 441 3375 450
rect 3339 439 3379 441
rect 3343 435 3345 439
rect 3349 435 3351 439
rect 3355 435 3357 439
rect 3361 435 3363 439
rect 3367 435 3369 439
rect 3373 435 3375 439
rect 3339 433 3379 435
rect 3343 429 3345 433
rect 3349 429 3351 433
rect 3355 429 3357 433
rect 3361 429 3363 433
rect 3367 429 3369 433
rect 3373 429 3375 433
rect 3339 427 3379 429
rect 3343 423 3345 427
rect 3349 423 3351 427
rect 3355 423 3357 427
rect 3361 423 3363 427
rect 3367 423 3369 427
rect 3373 423 3375 427
rect 3339 421 3379 423
rect 3343 412 3345 421
rect 3349 412 3351 421
rect 3355 412 3357 421
rect 3361 412 3363 421
rect 3367 412 3369 421
rect 3373 412 3375 421
rect 3387 509 3389 513
rect 3393 509 3395 513
rect 3399 509 3401 513
rect 3405 509 3407 513
rect 3411 509 3413 513
rect 3417 509 3419 513
rect 3383 499 3423 509
rect 3383 495 3389 499
rect 3393 495 3395 499
rect 3399 495 3401 499
rect 3405 495 3407 499
rect 3411 495 3413 499
rect 3417 495 3419 499
rect 3383 493 3423 495
rect 3387 489 3389 493
rect 3393 489 3395 493
rect 3399 489 3401 493
rect 3405 489 3407 493
rect 3411 489 3413 493
rect 3417 489 3419 493
rect 3383 487 3423 489
rect 3387 483 3389 487
rect 3393 483 3395 487
rect 3399 483 3401 487
rect 3405 483 3407 487
rect 3411 483 3413 487
rect 3417 483 3419 487
rect 3383 481 3423 483
rect 3387 477 3389 481
rect 3393 477 3395 481
rect 3399 477 3401 481
rect 3405 477 3407 481
rect 3411 477 3413 481
rect 3417 477 3419 481
rect 3383 475 3423 477
rect 3387 471 3389 475
rect 3393 471 3395 475
rect 3399 471 3401 475
rect 3405 471 3407 475
rect 3411 471 3413 475
rect 3417 471 3419 475
rect 3383 469 3423 471
rect 3387 465 3389 469
rect 3393 465 3395 469
rect 3399 465 3401 469
rect 3405 465 3407 469
rect 3411 465 3413 469
rect 3417 465 3419 469
rect 3383 449 3413 465
rect 3427 461 3436 509
rect 3417 460 3436 461
rect 3421 456 3422 460
rect 3426 456 3427 460
rect 3431 456 3432 460
rect 3417 455 3436 456
rect 3460 461 3469 509
rect 3477 509 3479 513
rect 3483 509 3485 513
rect 3489 509 3491 513
rect 3495 509 3497 513
rect 3501 509 3503 513
rect 3507 509 3509 513
rect 3473 499 3513 509
rect 3477 495 3479 499
rect 3483 495 3485 499
rect 3489 495 3491 499
rect 3495 495 3497 499
rect 3501 495 3503 499
rect 3507 495 3513 499
rect 3473 493 3513 495
rect 3477 489 3479 493
rect 3483 489 3485 493
rect 3489 489 3491 493
rect 3495 489 3497 493
rect 3501 489 3503 493
rect 3507 489 3509 493
rect 3473 487 3513 489
rect 3477 483 3479 487
rect 3483 483 3485 487
rect 3489 483 3491 487
rect 3495 483 3497 487
rect 3501 483 3503 487
rect 3507 483 3509 487
rect 3473 481 3513 483
rect 3477 477 3479 481
rect 3483 477 3485 481
rect 3489 477 3491 481
rect 3495 477 3497 481
rect 3501 477 3503 481
rect 3507 477 3509 481
rect 3473 475 3513 477
rect 3477 471 3479 475
rect 3483 471 3485 475
rect 3489 471 3491 475
rect 3495 471 3497 475
rect 3501 471 3503 475
rect 3507 471 3509 475
rect 3473 469 3513 471
rect 3477 465 3479 469
rect 3483 465 3485 469
rect 3489 465 3491 469
rect 3495 465 3497 469
rect 3501 465 3503 469
rect 3507 465 3509 469
rect 3460 460 3479 461
rect 3464 456 3465 460
rect 3469 456 3470 460
rect 3474 456 3475 460
rect 3460 455 3479 456
rect 3383 445 3384 449
rect 3388 445 3390 449
rect 3394 445 3396 449
rect 3400 445 3402 449
rect 3406 445 3408 449
rect 3412 445 3413 449
rect 3383 443 3413 445
rect 3383 439 3384 443
rect 3388 439 3390 443
rect 3394 439 3396 443
rect 3400 439 3402 443
rect 3406 439 3408 443
rect 3412 439 3413 443
rect 3383 437 3413 439
rect 3383 433 3384 437
rect 3388 433 3390 437
rect 3394 433 3396 437
rect 3400 433 3402 437
rect 3406 433 3408 437
rect 3412 433 3413 437
rect 3383 431 3413 433
rect 3383 427 3384 431
rect 3388 427 3390 431
rect 3394 427 3396 431
rect 3400 427 3402 431
rect 3406 427 3408 431
rect 3412 427 3413 431
rect 3383 424 3413 427
rect 3383 420 3384 424
rect 3388 420 3390 424
rect 3394 420 3396 424
rect 3400 420 3402 424
rect 3406 420 3408 424
rect 3412 420 3413 424
rect 3383 418 3413 420
rect 3383 414 3384 418
rect 3388 414 3390 418
rect 3394 414 3396 418
rect 3400 414 3402 418
rect 3406 414 3408 418
rect 3412 414 3413 418
rect 3383 413 3413 414
rect 3483 449 3513 465
rect 3483 445 3484 449
rect 3488 445 3490 449
rect 3494 445 3496 449
rect 3500 445 3502 449
rect 3506 445 3508 449
rect 3512 445 3513 449
rect 3483 443 3513 445
rect 3483 439 3484 443
rect 3488 439 3490 443
rect 3494 439 3496 443
rect 3500 439 3502 443
rect 3506 439 3508 443
rect 3512 439 3513 443
rect 3483 437 3513 439
rect 3483 433 3484 437
rect 3488 433 3490 437
rect 3494 433 3496 437
rect 3500 433 3502 437
rect 3506 433 3508 437
rect 3512 433 3513 437
rect 3483 431 3513 433
rect 3483 427 3484 431
rect 3488 427 3490 431
rect 3494 427 3496 431
rect 3500 427 3502 431
rect 3506 427 3508 431
rect 3512 427 3513 431
rect 3483 424 3513 427
rect 3483 420 3484 424
rect 3488 420 3490 424
rect 3494 420 3496 424
rect 3500 420 3502 424
rect 3506 420 3508 424
rect 3512 420 3513 424
rect 3483 418 3513 420
rect 3483 414 3484 418
rect 3488 414 3490 418
rect 3494 414 3496 418
rect 3500 414 3502 418
rect 3506 414 3508 418
rect 3512 414 3513 418
rect 3483 413 3513 414
rect 3521 509 3523 513
rect 3527 509 3529 513
rect 3533 509 3535 513
rect 3539 509 3541 513
rect 3545 509 3547 513
rect 3551 509 3553 513
rect 3517 505 3557 509
rect 3521 501 3523 505
rect 3527 501 3529 505
rect 3533 501 3535 505
rect 3539 501 3541 505
rect 3545 501 3547 505
rect 3551 501 3553 505
rect 3517 450 3557 501
rect 3521 441 3523 450
rect 3527 441 3529 450
rect 3533 441 3535 450
rect 3539 441 3541 450
rect 3545 441 3547 450
rect 3551 441 3553 450
rect 3517 439 3557 441
rect 3521 435 3523 439
rect 3527 435 3529 439
rect 3533 435 3535 439
rect 3539 435 3541 439
rect 3545 435 3547 439
rect 3551 435 3553 439
rect 3517 433 3557 435
rect 3521 429 3523 433
rect 3527 429 3529 433
rect 3533 429 3535 433
rect 3539 429 3541 433
rect 3545 429 3547 433
rect 3551 429 3553 433
rect 3517 427 3557 429
rect 3521 423 3523 427
rect 3527 423 3529 427
rect 3533 423 3535 427
rect 3539 423 3541 427
rect 3545 423 3547 427
rect 3551 423 3553 427
rect 3517 421 3557 423
rect 3339 376 3379 412
rect 3521 412 3523 421
rect 3527 412 3529 421
rect 3533 412 3535 421
rect 3539 412 3541 421
rect 3545 412 3547 421
rect 3551 412 3553 421
rect 3387 402 3389 406
rect 3393 402 3395 406
rect 3399 402 3401 406
rect 3405 402 3407 406
rect 3411 402 3413 406
rect 3417 402 3419 406
rect 3383 401 3423 402
rect 3387 397 3389 401
rect 3393 397 3395 401
rect 3399 397 3401 401
rect 3405 397 3407 401
rect 3411 397 3413 401
rect 3417 397 3419 401
rect 3383 394 3423 397
rect 3387 390 3389 394
rect 3393 390 3395 394
rect 3399 390 3401 394
rect 3405 390 3407 394
rect 3411 390 3413 394
rect 3417 390 3419 394
rect 3383 388 3423 390
rect 3387 384 3389 388
rect 3393 384 3395 388
rect 3399 384 3401 388
rect 3405 384 3407 388
rect 3411 384 3413 388
rect 3417 384 3419 388
rect 3389 382 3423 384
rect 3393 378 3395 382
rect 3399 378 3401 382
rect 3405 378 3407 382
rect 3411 378 3413 382
rect 3417 378 3419 382
rect 3477 402 3479 406
rect 3483 402 3485 406
rect 3489 402 3491 406
rect 3495 402 3497 406
rect 3501 402 3503 406
rect 3507 402 3509 406
rect 3473 401 3513 402
rect 3477 397 3479 401
rect 3483 397 3485 401
rect 3489 397 3491 401
rect 3495 397 3497 401
rect 3501 397 3503 401
rect 3507 397 3509 401
rect 3473 394 3513 397
rect 3477 390 3479 394
rect 3483 390 3485 394
rect 3489 390 3491 394
rect 3495 390 3497 394
rect 3501 390 3503 394
rect 3507 390 3509 394
rect 3473 388 3513 390
rect 3477 384 3479 388
rect 3483 384 3485 388
rect 3489 384 3491 388
rect 3495 384 3497 388
rect 3501 384 3503 388
rect 3507 384 3509 388
rect 3473 382 3507 384
rect 3477 378 3479 382
rect 3483 378 3485 382
rect 3489 378 3491 382
rect 3495 378 3497 382
rect 3501 378 3503 382
rect 3343 372 3345 376
rect 3349 372 3351 376
rect 3355 372 3357 376
rect 3361 372 3363 376
rect 3367 372 3369 376
rect 3373 372 3375 376
rect 3339 369 3379 372
rect 3517 376 3557 412
rect 3521 372 3523 376
rect 3527 372 3529 376
rect 3533 372 3535 376
rect 3539 372 3541 376
rect 3545 372 3547 376
rect 3551 372 3553 376
rect 3517 369 3557 372
rect 3817 509 3819 513
rect 3823 509 3825 513
rect 3829 509 3831 513
rect 3835 509 3837 513
rect 3841 509 3843 513
rect 3847 509 3849 513
rect 3813 505 3853 509
rect 3817 501 3819 505
rect 3823 501 3825 505
rect 3829 501 3831 505
rect 3835 501 3837 505
rect 3841 501 3843 505
rect 3847 501 3849 505
rect 3813 450 3853 501
rect 3817 441 3819 450
rect 3823 441 3825 450
rect 3829 441 3831 450
rect 3835 441 3837 450
rect 3841 441 3843 450
rect 3847 441 3849 450
rect 3813 439 3853 441
rect 3817 435 3819 439
rect 3823 435 3825 439
rect 3829 435 3831 439
rect 3835 435 3837 439
rect 3841 435 3843 439
rect 3847 435 3849 439
rect 3813 433 3853 435
rect 3817 429 3819 433
rect 3823 429 3825 433
rect 3829 429 3831 433
rect 3835 429 3837 433
rect 3841 429 3843 433
rect 3847 429 3849 433
rect 3813 427 3853 429
rect 3817 423 3819 427
rect 3823 423 3825 427
rect 3829 423 3831 427
rect 3835 423 3837 427
rect 3841 423 3843 427
rect 3847 423 3849 427
rect 3813 421 3853 423
rect 3817 412 3819 421
rect 3823 412 3825 421
rect 3829 412 3831 421
rect 3835 412 3837 421
rect 3841 412 3843 421
rect 3847 412 3849 421
rect 3861 509 3863 513
rect 3867 509 3869 513
rect 3873 509 3875 513
rect 3879 509 3881 513
rect 3885 509 3887 513
rect 3891 509 3893 513
rect 3857 499 3897 509
rect 3857 495 3863 499
rect 3867 495 3869 499
rect 3873 495 3875 499
rect 3879 495 3881 499
rect 3885 495 3887 499
rect 3891 495 3893 499
rect 3857 493 3897 495
rect 3861 489 3863 493
rect 3867 489 3869 493
rect 3873 489 3875 493
rect 3879 489 3881 493
rect 3885 489 3887 493
rect 3891 489 3893 493
rect 3857 487 3897 489
rect 3861 483 3863 487
rect 3867 483 3869 487
rect 3873 483 3875 487
rect 3879 483 3881 487
rect 3885 483 3887 487
rect 3891 483 3893 487
rect 3857 481 3897 483
rect 3861 477 3863 481
rect 3867 477 3869 481
rect 3873 477 3875 481
rect 3879 477 3881 481
rect 3885 477 3887 481
rect 3891 477 3893 481
rect 3857 475 3897 477
rect 3861 471 3863 475
rect 3867 471 3869 475
rect 3873 471 3875 475
rect 3879 471 3881 475
rect 3885 471 3887 475
rect 3891 471 3893 475
rect 3857 469 3897 471
rect 3861 465 3863 469
rect 3867 465 3869 469
rect 3873 465 3875 469
rect 3879 465 3881 469
rect 3885 465 3887 469
rect 3891 465 3893 469
rect 3857 449 3887 465
rect 3901 461 3910 509
rect 3891 460 3910 461
rect 3895 456 3896 460
rect 3900 456 3901 460
rect 3905 456 3906 460
rect 3891 455 3910 456
rect 3934 461 3943 509
rect 3951 509 3953 513
rect 3957 509 3959 513
rect 3963 509 3965 513
rect 3969 509 3971 513
rect 3975 509 3977 513
rect 3981 509 3983 513
rect 3947 499 3987 509
rect 3951 495 3953 499
rect 3957 495 3959 499
rect 3963 495 3965 499
rect 3969 495 3971 499
rect 3975 495 3977 499
rect 3981 495 3987 499
rect 3947 493 3987 495
rect 3951 489 3953 493
rect 3957 489 3959 493
rect 3963 489 3965 493
rect 3969 489 3971 493
rect 3975 489 3977 493
rect 3981 489 3983 493
rect 3947 487 3987 489
rect 3951 483 3953 487
rect 3957 483 3959 487
rect 3963 483 3965 487
rect 3969 483 3971 487
rect 3975 483 3977 487
rect 3981 483 3983 487
rect 3947 481 3987 483
rect 3951 477 3953 481
rect 3957 477 3959 481
rect 3963 477 3965 481
rect 3969 477 3971 481
rect 3975 477 3977 481
rect 3981 477 3983 481
rect 3947 475 3987 477
rect 3951 471 3953 475
rect 3957 471 3959 475
rect 3963 471 3965 475
rect 3969 471 3971 475
rect 3975 471 3977 475
rect 3981 471 3983 475
rect 3947 469 3987 471
rect 3951 465 3953 469
rect 3957 465 3959 469
rect 3963 465 3965 469
rect 3969 465 3971 469
rect 3975 465 3977 469
rect 3981 465 3983 469
rect 3934 460 3953 461
rect 3938 456 3939 460
rect 3943 456 3944 460
rect 3948 456 3949 460
rect 3934 455 3953 456
rect 3857 445 3858 449
rect 3862 445 3864 449
rect 3868 445 3870 449
rect 3874 445 3876 449
rect 3880 445 3882 449
rect 3886 445 3887 449
rect 3857 443 3887 445
rect 3857 439 3858 443
rect 3862 439 3864 443
rect 3868 439 3870 443
rect 3874 439 3876 443
rect 3880 439 3882 443
rect 3886 439 3887 443
rect 3857 437 3887 439
rect 3857 433 3858 437
rect 3862 433 3864 437
rect 3868 433 3870 437
rect 3874 433 3876 437
rect 3880 433 3882 437
rect 3886 433 3887 437
rect 3857 431 3887 433
rect 3857 427 3858 431
rect 3862 427 3864 431
rect 3868 427 3870 431
rect 3874 427 3876 431
rect 3880 427 3882 431
rect 3886 427 3887 431
rect 3857 424 3887 427
rect 3857 420 3858 424
rect 3862 420 3864 424
rect 3868 420 3870 424
rect 3874 420 3876 424
rect 3880 420 3882 424
rect 3886 420 3887 424
rect 3857 418 3887 420
rect 3857 414 3858 418
rect 3862 414 3864 418
rect 3868 414 3870 418
rect 3874 414 3876 418
rect 3880 414 3882 418
rect 3886 414 3887 418
rect 3857 413 3887 414
rect 3957 449 3987 465
rect 3957 445 3958 449
rect 3962 445 3964 449
rect 3968 445 3970 449
rect 3974 445 3976 449
rect 3980 445 3982 449
rect 3986 445 3987 449
rect 3957 443 3987 445
rect 3957 439 3958 443
rect 3962 439 3964 443
rect 3968 439 3970 443
rect 3974 439 3976 443
rect 3980 439 3982 443
rect 3986 439 3987 443
rect 3957 437 3987 439
rect 3957 433 3958 437
rect 3962 433 3964 437
rect 3968 433 3970 437
rect 3974 433 3976 437
rect 3980 433 3982 437
rect 3986 433 3987 437
rect 3957 431 3987 433
rect 3957 427 3958 431
rect 3962 427 3964 431
rect 3968 427 3970 431
rect 3974 427 3976 431
rect 3980 427 3982 431
rect 3986 427 3987 431
rect 3957 424 3987 427
rect 3957 420 3958 424
rect 3962 420 3964 424
rect 3968 420 3970 424
rect 3974 420 3976 424
rect 3980 420 3982 424
rect 3986 420 3987 424
rect 3957 418 3987 420
rect 3957 414 3958 418
rect 3962 414 3964 418
rect 3968 414 3970 418
rect 3974 414 3976 418
rect 3980 414 3982 418
rect 3986 414 3987 418
rect 3957 413 3987 414
rect 3995 509 3997 513
rect 4001 509 4003 513
rect 4007 509 4009 513
rect 4013 509 4015 513
rect 4019 509 4021 513
rect 4025 509 4027 513
rect 3991 505 4031 509
rect 3995 501 3997 505
rect 4001 501 4003 505
rect 4007 501 4009 505
rect 4013 501 4015 505
rect 4019 501 4021 505
rect 4025 501 4027 505
rect 3991 450 4031 501
rect 3995 441 3997 450
rect 4001 441 4003 450
rect 4007 441 4009 450
rect 4013 441 4015 450
rect 4019 441 4021 450
rect 4025 441 4027 450
rect 3991 439 4031 441
rect 3995 435 3997 439
rect 4001 435 4003 439
rect 4007 435 4009 439
rect 4013 435 4015 439
rect 4019 435 4021 439
rect 4025 435 4027 439
rect 3991 433 4031 435
rect 3995 429 3997 433
rect 4001 429 4003 433
rect 4007 429 4009 433
rect 4013 429 4015 433
rect 4019 429 4021 433
rect 4025 429 4027 433
rect 3991 427 4031 429
rect 3995 423 3997 427
rect 4001 423 4003 427
rect 4007 423 4009 427
rect 4013 423 4015 427
rect 4019 423 4021 427
rect 4025 423 4027 427
rect 3991 421 4031 423
rect 3813 376 3853 412
rect 3995 412 3997 421
rect 4001 412 4003 421
rect 4007 412 4009 421
rect 4013 412 4015 421
rect 4019 412 4021 421
rect 4025 412 4027 421
rect 3861 402 3863 406
rect 3867 402 3869 406
rect 3873 402 3875 406
rect 3879 402 3881 406
rect 3885 402 3887 406
rect 3891 402 3893 406
rect 3857 401 3897 402
rect 3861 397 3863 401
rect 3867 397 3869 401
rect 3873 397 3875 401
rect 3879 397 3881 401
rect 3885 397 3887 401
rect 3891 397 3893 401
rect 3857 394 3897 397
rect 3861 390 3863 394
rect 3867 390 3869 394
rect 3873 390 3875 394
rect 3879 390 3881 394
rect 3885 390 3887 394
rect 3891 390 3893 394
rect 3857 388 3897 390
rect 3861 384 3863 388
rect 3867 384 3869 388
rect 3873 384 3875 388
rect 3879 384 3881 388
rect 3885 384 3887 388
rect 3891 384 3893 388
rect 3863 382 3897 384
rect 3867 378 3869 382
rect 3873 378 3875 382
rect 3879 378 3881 382
rect 3885 378 3887 382
rect 3891 378 3893 382
rect 3951 402 3953 406
rect 3957 402 3959 406
rect 3963 402 3965 406
rect 3969 402 3971 406
rect 3975 402 3977 406
rect 3981 402 3983 406
rect 3947 401 3987 402
rect 3951 397 3953 401
rect 3957 397 3959 401
rect 3963 397 3965 401
rect 3969 397 3971 401
rect 3975 397 3977 401
rect 3981 397 3983 401
rect 3947 394 3987 397
rect 3951 390 3953 394
rect 3957 390 3959 394
rect 3963 390 3965 394
rect 3969 390 3971 394
rect 3975 390 3977 394
rect 3981 390 3983 394
rect 3947 388 3987 390
rect 3951 384 3953 388
rect 3957 384 3959 388
rect 3963 384 3965 388
rect 3969 384 3971 388
rect 3975 384 3977 388
rect 3981 384 3983 388
rect 3947 382 3981 384
rect 3951 378 3953 382
rect 3957 378 3959 382
rect 3963 378 3965 382
rect 3969 378 3971 382
rect 3975 378 3977 382
rect 3817 372 3819 376
rect 3823 372 3825 376
rect 3829 372 3831 376
rect 3835 372 3837 376
rect 3841 372 3843 376
rect 3847 372 3849 376
rect 3813 369 3853 372
rect 3991 376 4031 412
rect 3995 372 3997 376
rect 4001 372 4003 376
rect 4007 372 4009 376
rect 4013 372 4015 376
rect 4019 372 4021 376
rect 4025 372 4027 376
rect 3991 369 4031 372
rect 4291 509 4293 513
rect 4297 509 4299 513
rect 4303 509 4305 513
rect 4309 509 4311 513
rect 4315 509 4317 513
rect 4321 509 4323 513
rect 4287 505 4327 509
rect 4291 501 4293 505
rect 4297 501 4299 505
rect 4303 501 4305 505
rect 4309 501 4311 505
rect 4315 501 4317 505
rect 4321 501 4323 505
rect 4287 450 4327 501
rect 4291 441 4293 450
rect 4297 441 4299 450
rect 4303 441 4305 450
rect 4309 441 4311 450
rect 4315 441 4317 450
rect 4321 441 4323 450
rect 4287 439 4327 441
rect 4291 435 4293 439
rect 4297 435 4299 439
rect 4303 435 4305 439
rect 4309 435 4311 439
rect 4315 435 4317 439
rect 4321 435 4323 439
rect 4287 433 4327 435
rect 4291 429 4293 433
rect 4297 429 4299 433
rect 4303 429 4305 433
rect 4309 429 4311 433
rect 4315 429 4317 433
rect 4321 429 4323 433
rect 4287 427 4327 429
rect 4291 423 4293 427
rect 4297 423 4299 427
rect 4303 423 4305 427
rect 4309 423 4311 427
rect 4315 423 4317 427
rect 4321 423 4323 427
rect 4287 421 4327 423
rect 4291 412 4293 421
rect 4297 412 4299 421
rect 4303 412 4305 421
rect 4309 412 4311 421
rect 4315 412 4317 421
rect 4321 412 4323 421
rect 4335 509 4337 513
rect 4341 509 4343 513
rect 4347 509 4349 513
rect 4353 509 4355 513
rect 4359 509 4361 513
rect 4365 509 4367 513
rect 4331 499 4371 509
rect 4331 495 4337 499
rect 4341 495 4343 499
rect 4347 495 4349 499
rect 4353 495 4355 499
rect 4359 495 4361 499
rect 4365 495 4367 499
rect 4331 493 4371 495
rect 4335 489 4337 493
rect 4341 489 4343 493
rect 4347 489 4349 493
rect 4353 489 4355 493
rect 4359 489 4361 493
rect 4365 489 4367 493
rect 4331 487 4371 489
rect 4335 483 4337 487
rect 4341 483 4343 487
rect 4347 483 4349 487
rect 4353 483 4355 487
rect 4359 483 4361 487
rect 4365 483 4367 487
rect 4331 481 4371 483
rect 4335 477 4337 481
rect 4341 477 4343 481
rect 4347 477 4349 481
rect 4353 477 4355 481
rect 4359 477 4361 481
rect 4365 477 4367 481
rect 4331 475 4371 477
rect 4335 471 4337 475
rect 4341 471 4343 475
rect 4347 471 4349 475
rect 4353 471 4355 475
rect 4359 471 4361 475
rect 4365 471 4367 475
rect 4331 469 4371 471
rect 4335 465 4337 469
rect 4341 465 4343 469
rect 4347 465 4349 469
rect 4353 465 4355 469
rect 4359 465 4361 469
rect 4365 465 4367 469
rect 4331 449 4361 465
rect 4375 461 4384 509
rect 4365 460 4384 461
rect 4369 456 4370 460
rect 4374 456 4375 460
rect 4379 456 4380 460
rect 4365 455 4384 456
rect 4408 461 4417 509
rect 4425 509 4427 513
rect 4431 509 4433 513
rect 4437 509 4439 513
rect 4443 509 4445 513
rect 4449 509 4451 513
rect 4455 509 4457 513
rect 4421 499 4461 509
rect 4425 495 4427 499
rect 4431 495 4433 499
rect 4437 495 4439 499
rect 4443 495 4445 499
rect 4449 495 4451 499
rect 4455 495 4457 499
rect 4421 493 4461 495
rect 4425 489 4427 493
rect 4431 489 4433 493
rect 4437 489 4439 493
rect 4443 489 4445 493
rect 4449 489 4451 493
rect 4455 489 4457 493
rect 4421 487 4461 489
rect 4425 483 4427 487
rect 4431 483 4433 487
rect 4437 483 4439 487
rect 4443 483 4445 487
rect 4449 483 4451 487
rect 4455 483 4457 487
rect 4421 481 4461 483
rect 4425 477 4427 481
rect 4431 477 4433 481
rect 4437 477 4439 481
rect 4443 477 4445 481
rect 4449 477 4451 481
rect 4455 477 4457 481
rect 4421 475 4461 477
rect 4425 471 4427 475
rect 4431 471 4433 475
rect 4437 471 4439 475
rect 4443 471 4445 475
rect 4449 471 4451 475
rect 4455 471 4457 475
rect 4421 469 4461 471
rect 4425 465 4427 469
rect 4431 465 4433 469
rect 4437 465 4439 469
rect 4443 465 4445 469
rect 4449 465 4451 469
rect 4455 465 4457 469
rect 4408 460 4427 461
rect 4412 456 4413 460
rect 4417 456 4418 460
rect 4422 456 4423 460
rect 4408 455 4427 456
rect 4331 445 4332 449
rect 4336 445 4338 449
rect 4342 445 4344 449
rect 4348 445 4350 449
rect 4354 445 4356 449
rect 4360 445 4361 449
rect 4331 443 4361 445
rect 4331 439 4332 443
rect 4336 439 4338 443
rect 4342 439 4344 443
rect 4348 439 4350 443
rect 4354 439 4356 443
rect 4360 439 4361 443
rect 4331 437 4361 439
rect 4331 433 4332 437
rect 4336 433 4338 437
rect 4342 433 4344 437
rect 4348 433 4350 437
rect 4354 433 4356 437
rect 4360 433 4361 437
rect 4331 431 4361 433
rect 4331 427 4332 431
rect 4336 427 4338 431
rect 4342 427 4344 431
rect 4348 427 4350 431
rect 4354 427 4356 431
rect 4360 427 4361 431
rect 4331 424 4361 427
rect 4331 420 4332 424
rect 4336 420 4338 424
rect 4342 420 4344 424
rect 4348 420 4350 424
rect 4354 420 4356 424
rect 4360 420 4361 424
rect 4331 418 4361 420
rect 4331 414 4332 418
rect 4336 414 4338 418
rect 4342 414 4344 418
rect 4348 414 4350 418
rect 4354 414 4356 418
rect 4360 414 4361 418
rect 4331 413 4361 414
rect 4431 449 4461 465
rect 4431 445 4432 449
rect 4436 445 4438 449
rect 4442 445 4444 449
rect 4448 445 4450 449
rect 4454 445 4456 449
rect 4460 445 4461 449
rect 4431 443 4461 445
rect 4431 439 4432 443
rect 4436 439 4438 443
rect 4442 439 4444 443
rect 4448 439 4450 443
rect 4454 439 4456 443
rect 4460 439 4461 443
rect 4431 437 4461 439
rect 4431 433 4432 437
rect 4436 433 4438 437
rect 4442 433 4444 437
rect 4448 433 4450 437
rect 4454 433 4456 437
rect 4460 433 4461 437
rect 4431 431 4461 433
rect 4431 427 4432 431
rect 4436 427 4438 431
rect 4442 427 4444 431
rect 4448 427 4450 431
rect 4454 427 4456 431
rect 4460 427 4461 431
rect 4431 424 4461 427
rect 4431 420 4432 424
rect 4436 420 4438 424
rect 4442 420 4444 424
rect 4448 420 4450 424
rect 4454 420 4456 424
rect 4460 420 4461 424
rect 4431 418 4461 420
rect 4431 414 4432 418
rect 4436 414 4438 418
rect 4442 414 4444 418
rect 4448 414 4450 418
rect 4454 414 4456 418
rect 4460 414 4461 418
rect 4431 413 4461 414
rect 4465 450 4505 451
rect 4469 441 4471 450
rect 4475 441 4477 450
rect 4481 441 4483 450
rect 4487 441 4489 450
rect 4493 441 4495 450
rect 4499 441 4501 450
rect 4465 439 4505 441
rect 4469 435 4471 439
rect 4475 435 4477 439
rect 4481 435 4483 439
rect 4487 435 4489 439
rect 4493 435 4495 439
rect 4499 435 4501 439
rect 4465 433 4505 435
rect 4469 429 4471 433
rect 4475 429 4477 433
rect 4481 429 4483 433
rect 4487 429 4489 433
rect 4493 429 4495 433
rect 4499 429 4501 433
rect 4465 427 4505 429
rect 4469 423 4471 427
rect 4475 423 4477 427
rect 4481 423 4483 427
rect 4487 423 4489 427
rect 4493 423 4495 427
rect 4499 423 4501 427
rect 4465 421 4505 423
rect 4287 376 4327 412
rect 4469 412 4471 421
rect 4475 412 4477 421
rect 4481 412 4483 421
rect 4487 412 4489 421
rect 4493 412 4495 421
rect 4499 412 4501 421
rect 4335 402 4337 406
rect 4341 402 4343 406
rect 4347 402 4349 406
rect 4353 402 4355 406
rect 4359 402 4361 406
rect 4365 402 4367 406
rect 4331 401 4371 402
rect 4335 397 4337 401
rect 4341 397 4343 401
rect 4347 397 4349 401
rect 4353 397 4355 401
rect 4359 397 4361 401
rect 4365 397 4367 401
rect 4331 394 4371 397
rect 4335 390 4337 394
rect 4341 390 4343 394
rect 4347 390 4349 394
rect 4353 390 4355 394
rect 4359 390 4361 394
rect 4365 390 4367 394
rect 4331 388 4371 390
rect 4335 384 4337 388
rect 4341 384 4343 388
rect 4347 384 4349 388
rect 4353 384 4355 388
rect 4359 384 4361 388
rect 4365 384 4367 388
rect 4337 382 4371 384
rect 4341 378 4343 382
rect 4347 378 4349 382
rect 4353 378 4355 382
rect 4359 378 4361 382
rect 4365 378 4367 382
rect 4425 402 4427 406
rect 4431 402 4433 406
rect 4437 402 4439 406
rect 4443 402 4445 406
rect 4449 402 4451 406
rect 4455 402 4457 406
rect 4421 401 4461 402
rect 4425 397 4427 401
rect 4431 397 4433 401
rect 4437 397 4439 401
rect 4443 397 4445 401
rect 4449 397 4451 401
rect 4455 397 4457 401
rect 4421 394 4461 397
rect 4425 390 4427 394
rect 4431 390 4433 394
rect 4437 390 4439 394
rect 4443 390 4445 394
rect 4449 390 4451 394
rect 4455 390 4457 394
rect 4421 388 4461 390
rect 4425 384 4427 388
rect 4431 384 4433 388
rect 4437 384 4439 388
rect 4443 384 4445 388
rect 4449 384 4451 388
rect 4455 384 4457 388
rect 4421 382 4455 384
rect 4425 378 4427 382
rect 4431 378 4433 382
rect 4437 378 4439 382
rect 4443 378 4445 382
rect 4449 378 4451 382
rect 4291 372 4293 376
rect 4297 372 4299 376
rect 4303 372 4305 376
rect 4309 372 4311 376
rect 4315 372 4317 376
rect 4321 372 4323 376
rect 4287 369 4327 372
rect 4465 376 4505 412
rect 4469 372 4471 376
rect 4475 372 4477 376
rect 4481 372 4483 376
rect 4487 372 4489 376
rect 4493 372 4495 376
rect 4499 372 4501 376
rect 4465 369 4505 372
rect 3 365 5 369
rect 9 365 11 369
rect 15 365 17 369
rect 21 365 23 369
rect 27 365 29 369
rect 33 365 35 369
rect 39 365 41 369
rect 45 365 47 369
rect 51 365 53 369
rect 57 365 59 369
rect 63 365 65 369
rect 69 365 71 369
rect 75 365 77 369
rect 81 365 83 369
rect 87 365 89 369
rect 93 365 95 369
rect 99 365 101 369
rect 105 365 107 369
rect 111 365 113 369
rect 117 365 119 369
rect 123 365 125 369
rect 129 365 131 369
rect 135 365 137 369
rect 141 365 143 369
rect 147 365 149 369
rect 153 365 155 369
rect 159 365 161 369
rect 165 365 167 369
rect 171 365 173 369
rect 177 365 179 369
rect 183 365 185 369
rect 189 365 191 369
rect 195 365 197 369
rect 201 365 203 369
rect 207 365 209 369
rect 213 365 215 369
rect 219 365 221 369
rect 225 365 227 369
rect 231 365 233 369
rect 237 365 239 369
rect 243 365 245 369
rect 249 365 251 369
rect 255 365 257 369
rect 261 365 263 369
rect 267 365 269 369
rect 273 365 275 369
rect 279 365 281 369
rect 285 365 287 369
rect 291 365 293 369
rect 297 365 299 369
rect 303 365 305 369
rect 309 365 311 369
rect 315 365 317 369
rect 321 365 323 369
rect 327 365 329 369
rect 333 365 335 369
rect 339 365 341 369
rect 345 365 347 369
rect 351 365 353 369
rect 357 365 359 369
rect 363 365 365 369
rect 369 365 371 369
rect 375 365 377 369
rect 381 365 383 369
rect 387 365 389 369
rect 393 365 395 369
rect 399 365 401 369
rect 405 365 407 369
rect 411 365 413 369
rect 417 365 419 369
rect 423 365 425 369
rect 429 365 431 369
rect 435 365 437 369
rect 441 365 443 369
rect 447 365 449 369
rect 453 365 455 369
rect 459 365 461 369
rect 465 365 467 369
rect 471 365 473 369
rect 477 365 479 369
rect 483 365 485 369
rect 489 365 491 369
rect 495 365 497 369
rect 501 365 503 369
rect 507 365 509 369
rect 513 365 515 369
rect 519 365 521 369
rect 525 365 527 369
rect 531 365 533 369
rect 537 365 539 369
rect 543 365 545 369
rect 549 365 551 369
rect 555 365 557 369
rect 561 365 563 369
rect 567 365 569 369
rect 573 365 575 369
rect 579 365 581 369
rect 585 365 587 369
rect 621 365 623 369
rect 627 365 629 369
rect 633 365 635 369
rect 639 365 641 369
rect 645 365 647 369
rect 651 365 653 369
rect 657 365 659 369
rect 663 365 665 369
rect 669 365 671 369
rect 675 365 677 369
rect 681 365 683 369
rect 687 365 689 369
rect 693 365 695 369
rect 699 365 701 369
rect 705 365 707 369
rect 711 365 713 369
rect 717 365 719 369
rect 723 365 725 369
rect 729 365 731 369
rect 735 365 737 369
rect 741 365 743 369
rect 747 365 749 369
rect 753 365 755 369
rect 759 365 761 369
rect 765 365 767 369
rect 771 365 773 369
rect 777 365 779 369
rect 783 365 785 369
rect 789 365 791 369
rect 795 365 797 369
rect 801 365 803 369
rect 807 365 809 369
rect 813 365 815 369
rect 819 365 821 369
rect 825 365 827 369
rect 831 365 833 369
rect 837 365 839 369
rect 843 365 845 369
rect 849 365 851 369
rect 855 365 857 369
rect 861 365 863 369
rect 867 365 869 369
rect 873 365 875 369
rect 879 365 881 369
rect 885 365 887 369
rect 891 365 893 369
rect 897 365 899 369
rect 903 365 905 369
rect 909 365 911 369
rect 915 365 917 369
rect 921 365 923 369
rect 927 365 929 369
rect 933 365 935 369
rect 939 365 941 369
rect 945 365 947 369
rect 951 365 953 369
rect 957 365 959 369
rect 963 365 965 369
rect 969 365 971 369
rect 975 365 977 369
rect 981 365 983 369
rect 987 365 989 369
rect 993 365 995 369
rect 999 365 1001 369
rect 1005 365 1007 369
rect 1011 365 1013 369
rect 1017 365 1019 369
rect 1023 365 1025 369
rect 1029 365 1031 369
rect 1035 365 1037 369
rect 1041 365 1043 369
rect 1047 365 1049 369
rect 1053 365 1055 369
rect 1059 365 1061 369
rect 1095 365 1097 369
rect 1101 365 1103 369
rect 1107 365 1109 369
rect 1113 365 1115 369
rect 1119 365 1121 369
rect 1125 365 1127 369
rect 1131 365 1133 369
rect 1137 365 1139 369
rect 1143 365 1145 369
rect 1149 365 1151 369
rect 1155 365 1157 369
rect 1161 365 1163 369
rect 1167 365 1169 369
rect 1173 365 1175 369
rect 1179 365 1181 369
rect 1185 365 1187 369
rect 1191 365 1193 369
rect 1197 365 1199 369
rect 1203 365 1205 369
rect 1209 365 1211 369
rect 1215 365 1217 369
rect 1221 365 1223 369
rect 1227 365 1229 369
rect 1233 365 1235 369
rect 1239 365 1241 369
rect 1245 365 1247 369
rect 1251 365 1253 369
rect 1257 365 1259 369
rect 1263 365 1265 369
rect 1269 365 1271 369
rect 1275 365 1277 369
rect 1281 365 1283 369
rect 1287 365 1289 369
rect 1293 365 1295 369
rect 1299 365 1301 369
rect 1305 365 1307 369
rect 1311 365 1313 369
rect 1317 365 1319 369
rect 1323 365 1325 369
rect 1329 365 1331 369
rect 1335 365 1337 369
rect 1341 365 1343 369
rect 1347 365 1349 369
rect 1353 365 1355 369
rect 1359 365 1361 369
rect 1365 365 1367 369
rect 1371 365 1373 369
rect 1377 365 1379 369
rect 1383 365 1385 369
rect 1389 365 1391 369
rect 1395 365 1397 369
rect 1401 365 1403 369
rect 1407 365 1409 369
rect 1413 365 1415 369
rect 1419 365 1421 369
rect 1425 365 1427 369
rect 1431 365 1433 369
rect 1437 365 1439 369
rect 1443 365 1445 369
rect 1449 365 1451 369
rect 1455 365 1457 369
rect 1461 365 1463 369
rect 1467 365 1469 369
rect 1473 365 1475 369
rect 1479 365 1481 369
rect 1485 365 1487 369
rect 1491 365 1493 369
rect 1497 365 1499 369
rect 1503 365 1505 369
rect 1509 365 1511 369
rect 1515 365 1517 369
rect 1521 365 1523 369
rect 1527 365 1529 369
rect 1533 365 1535 369
rect 1569 365 1571 369
rect 1575 365 1577 369
rect 1581 365 1583 369
rect 1587 365 1589 369
rect 1593 365 1595 369
rect 1599 365 1601 369
rect 1605 365 1607 369
rect 1611 365 1613 369
rect 1617 365 1619 369
rect 1623 365 1625 369
rect 1629 365 1631 369
rect 1635 365 1637 369
rect 1641 365 1643 369
rect 1647 365 1649 369
rect 1653 365 1655 369
rect 1659 365 1661 369
rect 1665 365 1667 369
rect 1671 365 1673 369
rect 1677 365 1679 369
rect 1683 365 1685 369
rect 1689 365 1691 369
rect 1695 365 1697 369
rect 1701 365 1703 369
rect 1707 365 1709 369
rect 1713 365 1715 369
rect 1719 365 1721 369
rect 1725 365 1727 369
rect 1731 365 1733 369
rect 1737 365 1739 369
rect 1743 365 1745 369
rect 1749 365 1751 369
rect 1755 365 1757 369
rect 1761 365 1763 369
rect 1767 365 1769 369
rect 1773 365 1775 369
rect 1779 365 1781 369
rect 1785 365 1787 369
rect 1791 365 1793 369
rect 1797 365 1799 369
rect 1803 365 1805 369
rect 1809 365 1811 369
rect 1815 365 1817 369
rect 1821 365 1823 369
rect 1827 365 1829 369
rect 1833 365 1835 369
rect 1839 365 1841 369
rect 1845 365 1847 369
rect 1851 365 1853 369
rect 1857 365 1859 369
rect 1863 365 1865 369
rect 1869 365 1871 369
rect 1875 365 1877 369
rect 1881 365 1883 369
rect 1887 365 1889 369
rect 1893 365 1895 369
rect 1899 365 1901 369
rect 1905 365 1907 369
rect 1911 365 1913 369
rect 1917 365 1919 369
rect 1923 365 1925 369
rect 1929 365 1931 369
rect 1935 365 1937 369
rect 1941 365 1943 369
rect 1947 365 1949 369
rect 1953 365 1955 369
rect 1959 365 1961 369
rect 1965 365 1967 369
rect 1971 365 1973 369
rect 1977 365 1979 369
rect 1983 365 1985 369
rect 1989 365 1991 369
rect 1995 365 1997 369
rect 2001 365 2003 369
rect 2007 365 2009 369
rect 2043 365 2045 369
rect 2049 365 2051 369
rect 2055 365 2057 369
rect 2061 365 2063 369
rect 2067 365 2069 369
rect 2073 365 2075 369
rect 2079 365 2081 369
rect 2085 365 2087 369
rect 2091 365 2093 369
rect 2097 365 2099 369
rect 2103 365 2105 369
rect 2109 365 2111 369
rect 2115 365 2117 369
rect 2121 365 2123 369
rect 2127 365 2129 369
rect 2133 365 2135 369
rect 2139 365 2141 369
rect 2145 365 2147 369
rect 2151 365 2153 369
rect 2157 365 2159 369
rect 2163 365 2165 369
rect 2169 365 2171 369
rect 2175 365 2177 369
rect 2181 365 2183 369
rect 2187 365 2189 369
rect 2193 365 2195 369
rect 2199 365 2201 369
rect 2205 365 2207 369
rect 2211 365 2213 369
rect 2217 365 2219 369
rect 2223 365 2225 369
rect 2229 365 2231 369
rect 2235 365 2237 369
rect 2241 365 2243 369
rect 2247 365 2249 369
rect 2253 365 2255 369
rect 2259 365 2261 369
rect 2265 365 2267 369
rect 2271 365 2273 369
rect 2277 365 2279 369
rect 2283 365 2285 369
rect 2289 365 2291 369
rect 2295 365 2297 369
rect 2301 365 2303 369
rect 2307 365 2309 369
rect 2313 365 2315 369
rect 2319 365 2321 369
rect 2325 365 2327 369
rect 2331 365 2333 369
rect 2337 365 2339 369
rect 2343 365 2345 369
rect 2349 365 2351 369
rect 2355 365 2357 369
rect 2361 365 2363 369
rect 2367 365 2369 369
rect 2373 365 2375 369
rect 2379 365 2381 369
rect 2385 365 2387 369
rect 2391 365 2393 369
rect 2397 365 2399 369
rect 2403 365 2405 369
rect 2409 365 2411 369
rect 2415 365 2417 369
rect 2421 365 2423 369
rect 2427 365 2429 369
rect 2433 365 2435 369
rect 2439 365 2441 369
rect 2445 365 2447 369
rect 2451 365 2453 369
rect 2457 365 2459 369
rect 2463 365 2465 369
rect 2469 365 2471 369
rect 2475 365 2477 369
rect 2481 365 2483 369
rect 2517 365 2519 369
rect 2523 365 2525 369
rect 2529 365 2531 369
rect 2535 365 2537 369
rect 2541 365 2543 369
rect 2547 365 2549 369
rect 2553 365 2555 369
rect 2559 365 2561 369
rect 2565 365 2567 369
rect 2571 365 2573 369
rect 2577 365 2579 369
rect 2583 365 2585 369
rect 2589 365 2591 369
rect 2595 365 2597 369
rect 2601 365 2603 369
rect 2607 365 2609 369
rect 2613 365 2615 369
rect 2619 365 2621 369
rect 2625 365 2627 369
rect 2631 365 2633 369
rect 2637 365 2639 369
rect 2643 365 2645 369
rect 2649 365 2651 369
rect 2655 365 2657 369
rect 2661 365 2663 369
rect 2667 365 2669 369
rect 2673 365 2675 369
rect 2679 365 2681 369
rect 2685 365 2687 369
rect 2691 365 2693 369
rect 2697 365 2699 369
rect 2703 365 2705 369
rect 2709 365 2711 369
rect 2715 365 2717 369
rect 2721 365 2723 369
rect 2727 365 2729 369
rect 2733 365 2735 369
rect 2739 365 2741 369
rect 2745 365 2747 369
rect 2751 365 2753 369
rect 2757 365 2759 369
rect 2763 365 2765 369
rect 2769 365 2771 369
rect 2775 365 2777 369
rect 2781 365 2783 369
rect 2787 365 2789 369
rect 2793 365 2795 369
rect 2799 365 2801 369
rect 2805 365 2807 369
rect 2811 365 2813 369
rect 2817 365 2819 369
rect 2823 365 2825 369
rect 2829 365 2831 369
rect 2835 365 2837 369
rect 2841 365 2843 369
rect 2847 365 2849 369
rect 2853 365 2855 369
rect 2859 365 2861 369
rect 2865 365 2867 369
rect 2871 365 2873 369
rect 2877 365 2879 369
rect 2883 365 2885 369
rect 2889 365 2891 369
rect 2895 365 2897 369
rect 2901 365 2903 369
rect 2907 365 2909 369
rect 2913 365 2915 369
rect 2919 365 2921 369
rect 2925 365 2927 369
rect 2931 365 2933 369
rect 2937 365 2939 369
rect 2943 365 2945 369
rect 2949 365 2951 369
rect 2955 365 2957 369
rect 2991 365 2993 369
rect 2997 365 2999 369
rect 3003 365 3005 369
rect 3009 365 3011 369
rect 3015 365 3017 369
rect 3021 365 3023 369
rect 3027 365 3029 369
rect 3033 365 3035 369
rect 3039 365 3041 369
rect 3045 365 3047 369
rect 3051 365 3053 369
rect 3057 365 3059 369
rect 3063 365 3065 369
rect 3069 365 3071 369
rect 3075 365 3077 369
rect 3081 365 3083 369
rect 3087 365 3089 369
rect 3093 365 3095 369
rect 3099 365 3101 369
rect 3105 365 3107 369
rect 3111 365 3113 369
rect 3117 365 3119 369
rect 3123 365 3125 369
rect 3129 365 3131 369
rect 3135 365 3137 369
rect 3141 365 3143 369
rect 3147 365 3149 369
rect 3153 365 3155 369
rect 3159 365 3161 369
rect 3165 365 3167 369
rect 3171 365 3173 369
rect 3177 365 3179 369
rect 3183 365 3185 369
rect 3189 365 3191 369
rect 3195 365 3197 369
rect 3201 365 3203 369
rect 3207 365 3209 369
rect 3213 365 3215 369
rect 3219 365 3221 369
rect 3225 365 3227 369
rect 3231 365 3233 369
rect 3237 365 3239 369
rect 3243 365 3245 369
rect 3249 365 3251 369
rect 3255 365 3257 369
rect 3261 365 3263 369
rect 3267 365 3269 369
rect 3273 365 3275 369
rect 3279 365 3281 369
rect 3285 365 3287 369
rect 3291 365 3293 369
rect 3297 365 3299 369
rect 3303 365 3305 369
rect 3309 365 3311 369
rect 3315 365 3317 369
rect 3321 365 3323 369
rect 3327 365 3329 369
rect 3333 365 3335 369
rect 3339 365 3341 369
rect 3345 365 3347 369
rect 3351 365 3353 369
rect 3357 365 3359 369
rect 3363 365 3365 369
rect 3369 365 3371 369
rect 3375 365 3377 369
rect 3381 365 3383 369
rect 3387 365 3389 369
rect 3393 365 3395 369
rect 3399 365 3401 369
rect 3405 365 3407 369
rect 3411 365 3413 369
rect 3417 365 3419 369
rect 3423 365 3425 369
rect 3429 365 3431 369
rect 3465 365 3467 369
rect 3471 365 3473 369
rect 3477 365 3479 369
rect 3483 365 3485 369
rect 3489 365 3491 369
rect 3495 365 3497 369
rect 3501 365 3503 369
rect 3507 365 3509 369
rect 3513 365 3515 369
rect 3519 365 3521 369
rect 3525 365 3527 369
rect 3531 365 3533 369
rect 3537 365 3539 369
rect 3543 365 3545 369
rect 3549 365 3551 369
rect 3555 365 3557 369
rect 3561 365 3563 369
rect 3567 365 3569 369
rect 3573 365 3575 369
rect 3579 365 3581 369
rect 3585 365 3587 369
rect 3591 365 3593 369
rect 3597 365 3599 369
rect 3603 365 3605 369
rect 3609 365 3611 369
rect 3615 365 3617 369
rect 3621 365 3623 369
rect 3627 365 3629 369
rect 3633 365 3635 369
rect 3639 365 3641 369
rect 3645 365 3647 369
rect 3651 365 3653 369
rect 3657 365 3659 369
rect 3663 365 3665 369
rect 3669 365 3671 369
rect 3675 365 3677 369
rect 3681 365 3683 369
rect 3687 365 3689 369
rect 3693 365 3695 369
rect 3699 365 3701 369
rect 3705 365 3707 369
rect 3711 365 3713 369
rect 3717 365 3719 369
rect 3723 365 3725 369
rect 3729 365 3731 369
rect 3735 365 3737 369
rect 3741 365 3743 369
rect 3747 365 3749 369
rect 3753 365 3755 369
rect 3759 365 3761 369
rect 3765 365 3767 369
rect 3771 365 3773 369
rect 3777 365 3779 369
rect 3783 365 3785 369
rect 3789 365 3791 369
rect 3795 365 3797 369
rect 3801 365 3803 369
rect 3807 365 3809 369
rect 3813 365 3815 369
rect 3819 365 3821 369
rect 3825 365 3827 369
rect 3831 365 3833 369
rect 3837 365 3839 369
rect 3843 365 3845 369
rect 3849 365 3851 369
rect 3855 365 3857 369
rect 3861 365 3863 369
rect 3867 365 3869 369
rect 3873 365 3875 369
rect 3879 365 3881 369
rect 3885 365 3887 369
rect 3891 365 3893 369
rect 3897 365 3899 369
rect 3903 365 3905 369
rect 3939 365 3941 369
rect 3945 365 3947 369
rect 3951 365 3953 369
rect 3957 365 3959 369
rect 3963 365 3965 369
rect 3969 365 3971 369
rect 3975 365 3977 369
rect 3981 365 3983 369
rect 3987 365 3989 369
rect 3993 365 3995 369
rect 3999 365 4001 369
rect 4005 365 4007 369
rect 4011 365 4013 369
rect 4017 365 4019 369
rect 4023 365 4025 369
rect 4029 365 4031 369
rect 4035 365 4037 369
rect 4041 365 4043 369
rect 4047 365 4049 369
rect 4053 365 4055 369
rect 4059 365 4061 369
rect 4065 365 4067 369
rect 4071 365 4073 369
rect 4077 365 4079 369
rect 4083 365 4085 369
rect 4089 365 4091 369
rect 4095 365 4097 369
rect 4101 365 4103 369
rect 4107 365 4109 369
rect 4113 365 4115 369
rect 4119 365 4121 369
rect 4125 365 4127 369
rect 4131 365 4133 369
rect 4137 365 4139 369
rect 4143 365 4145 369
rect 4149 365 4151 369
rect 4155 365 4157 369
rect 4161 365 4163 369
rect 4167 365 4169 369
rect 4173 365 4175 369
rect 4179 365 4181 369
rect 4185 365 4187 369
rect 4191 365 4193 369
rect 4197 365 4199 369
rect 4203 365 4205 369
rect 4209 365 4211 369
rect 4215 365 4217 369
rect 4221 365 4223 369
rect 4227 365 4229 369
rect 4233 365 4235 369
rect 4239 365 4241 369
rect 4245 365 4247 369
rect 4251 365 4253 369
rect 4257 365 4259 369
rect 4263 365 4265 369
rect 4269 365 4271 369
rect 4275 365 4277 369
rect 4281 365 4283 369
rect 4287 365 4289 369
rect 4293 365 4295 369
rect 4299 365 4301 369
rect 4305 365 4307 369
rect 4311 365 4313 369
rect 4317 365 4319 369
rect 4323 365 4325 369
rect 4329 365 4331 369
rect 4335 365 4337 369
rect 4341 365 4343 369
rect 4347 365 4349 369
rect 4353 365 4355 369
rect 4359 365 4361 369
rect 4365 365 4367 369
rect 4371 365 4373 369
rect 4377 365 4379 369
rect 4413 365 4415 369
rect 4419 365 4421 369
rect 4425 365 4427 369
rect 4431 365 4433 369
rect 4437 365 4439 369
rect 4443 365 4445 369
rect 4449 365 4451 369
rect 4455 365 4457 369
rect 4461 365 4463 369
rect 4467 365 4469 369
rect 4473 365 4475 369
rect 4479 365 4481 369
rect 4485 365 4487 369
rect 4491 365 4493 369
rect 4497 365 4499 369
rect 4503 365 4505 369
rect 4509 365 4511 369
rect 4515 365 4517 369
rect 4521 365 4523 369
rect 4527 365 4529 369
rect 4533 365 4535 369
rect 4539 365 4541 369
rect 4545 365 4547 369
rect 4551 365 4553 369
rect 4557 365 4559 369
rect 4563 365 4565 369
rect 4569 365 4571 369
rect 4575 365 4577 369
rect 4581 365 4583 369
rect 4587 365 4589 369
rect 4593 365 4595 369
rect 4599 365 4601 369
rect 4605 365 4607 369
rect 4611 365 4613 369
rect 4617 365 4619 369
rect 4623 365 4625 369
rect 4629 365 4631 369
rect 4635 365 4637 369
rect 4641 365 4643 369
rect 4647 365 4649 369
rect 4653 365 4655 369
rect 4659 365 4661 369
rect 4665 365 4667 369
rect 4671 365 4673 369
rect 4677 365 4679 369
rect 4683 365 4685 369
rect 4689 365 4691 369
rect 4695 365 4697 369
rect 4701 365 4703 369
rect 4707 365 4709 369
rect 4713 365 4715 369
rect 4719 365 4721 369
rect 4725 365 4727 369
rect 4731 365 4733 369
rect 4737 365 4739 369
rect 4743 365 4745 369
rect 4749 365 4751 369
rect 4755 365 4757 369
rect 4761 365 4763 369
rect 4767 365 4769 369
rect 4773 365 4775 369
rect 4779 365 4781 369
rect 4785 365 4787 369
rect 4791 365 4793 369
rect 4797 365 4799 369
rect 4803 365 4805 369
rect 4809 365 4811 369
rect 4815 365 4817 369
rect 4821 365 4823 369
rect 4827 365 4829 369
rect 4833 365 4835 369
rect 4839 365 4841 369
rect 4845 365 4847 369
rect 4851 365 4853 369
rect 4857 365 4859 369
rect 4863 365 4865 369
rect 4869 365 4871 369
rect 4875 365 4877 369
rect 4881 365 4883 369
rect 4887 365 4889 369
rect 4893 365 4895 369
rect 4899 365 4901 369
rect 4905 365 4907 369
rect 4911 365 4913 369
rect 4917 365 4919 369
rect 4923 365 4925 369
rect 4929 365 4931 369
rect 4935 365 4937 369
rect 4941 365 4943 369
rect 4947 365 4949 369
rect 4953 365 4955 369
rect 4959 365 4961 369
rect 4965 365 4967 369
rect 4971 365 4973 369
rect 4977 365 4979 369
rect 4983 365 4985 369
rect 4989 365 4991 369
rect 4995 365 4997 369
rect 3 362 7 365
rect 323 363 369 365
rect 323 362 365 363
rect 327 358 329 362
rect 333 358 335 362
rect 339 358 341 362
rect 345 358 347 362
rect 351 358 353 362
rect 357 359 365 362
rect 357 358 369 359
rect 3 356 7 358
rect 3 350 7 352
rect 3 344 7 346
rect 3 338 7 340
rect 3 332 7 334
rect 3 326 7 328
rect 358 357 369 358
rect 362 353 365 357
rect 358 351 369 353
rect 362 347 365 351
rect 358 345 369 347
rect 362 341 365 345
rect 358 339 369 341
rect 362 335 365 339
rect 358 333 369 335
rect 362 329 365 333
rect 358 327 369 329
rect 362 323 365 327
rect 3 320 7 322
rect 365 321 369 323
rect 365 315 369 317
rect 365 309 369 311
rect 365 303 369 305
rect 365 297 369 299
rect 365 291 369 293
rect 365 285 369 287
rect 365 279 369 281
rect 365 273 369 275
rect 365 267 369 269
rect 365 261 369 263
rect 320 259 356 260
rect 320 255 327 259
rect 331 255 339 259
rect 343 255 351 259
rect 355 255 356 259
rect 320 253 356 255
rect 320 249 321 253
rect 325 249 327 253
rect 331 249 333 253
rect 337 249 339 253
rect 343 249 345 253
rect 349 249 351 253
rect 355 249 356 253
rect 320 247 356 249
rect 320 243 321 247
rect 325 243 333 247
rect 337 243 345 247
rect 349 243 356 247
rect 320 241 356 243
rect 320 237 321 241
rect 325 237 327 241
rect 331 237 333 241
rect 337 237 339 241
rect 343 237 345 241
rect 349 237 351 241
rect 355 237 356 241
rect 320 235 356 237
rect 320 231 327 235
rect 331 231 339 235
rect 343 231 351 235
rect 355 231 356 235
rect 320 229 356 231
rect 320 225 321 229
rect 325 225 327 229
rect 331 225 333 229
rect 337 225 339 229
rect 343 225 345 229
rect 349 225 351 229
rect 355 225 356 229
rect 320 223 356 225
rect 320 219 321 223
rect 325 219 333 223
rect 337 219 345 223
rect 349 219 356 223
rect 320 218 356 219
rect 365 255 369 257
rect 365 249 369 251
rect 365 243 369 245
rect 365 237 369 239
rect 365 231 369 233
rect 365 225 369 227
rect 365 219 369 221
rect 365 213 369 215
rect 365 207 369 209
rect 365 201 369 203
rect 365 195 369 197
rect 365 189 369 191
rect 365 183 369 185
rect 365 177 369 179
rect 365 171 369 173
rect 365 165 369 167
rect 365 159 369 161
rect 365 153 369 155
rect 365 147 369 149
rect 365 141 369 143
rect 365 135 369 137
rect 365 129 369 131
rect 365 123 369 125
rect 365 117 369 119
rect 365 111 369 113
rect 365 105 369 107
rect 365 99 369 101
rect 365 93 369 95
rect 365 87 369 89
rect 365 81 369 83
rect 365 75 369 77
rect 365 69 369 71
rect 365 63 369 65
rect 365 57 369 59
rect 365 51 369 53
rect 365 45 369 47
rect 365 39 369 41
rect 365 33 369 35
rect 365 27 369 29
rect 365 21 369 23
rect 365 15 369 17
rect 365 9 369 11
rect 320 3 322 7
rect 326 3 328 7
rect 332 3 334 7
rect 338 3 340 7
rect 344 3 346 7
rect 350 3 352 7
rect 356 3 358 7
rect 362 5 365 7
rect 362 3 369 5
rect 839 363 843 365
rect 839 357 843 359
rect 839 351 843 353
rect 839 345 843 347
rect 839 339 843 341
rect 839 333 843 335
rect 839 327 843 329
rect 839 321 843 323
rect 839 315 843 317
rect 839 309 843 311
rect 839 303 843 305
rect 839 297 843 299
rect 839 291 843 293
rect 839 285 843 287
rect 839 279 843 281
rect 839 273 843 275
rect 839 267 843 269
rect 839 261 843 263
rect 839 255 843 257
rect 839 249 843 251
rect 839 243 843 245
rect 839 237 843 239
rect 839 231 843 233
rect 839 225 843 227
rect 839 219 843 221
rect 839 213 843 215
rect 839 207 843 209
rect 839 201 843 203
rect 839 195 843 197
rect 839 189 843 191
rect 839 183 843 185
rect 839 177 843 179
rect 839 171 843 173
rect 839 165 843 167
rect 839 159 843 161
rect 839 153 843 155
rect 839 147 843 149
rect 839 141 843 143
rect 839 135 843 137
rect 839 129 843 131
rect 839 123 843 125
rect 839 117 843 119
rect 839 111 843 113
rect 839 105 843 107
rect 839 99 843 101
rect 839 93 843 95
rect 839 87 843 89
rect 839 81 843 83
rect 839 75 843 77
rect 839 69 843 71
rect 839 63 843 65
rect 839 57 843 59
rect 839 51 843 53
rect 839 45 843 47
rect 839 39 843 41
rect 839 33 843 35
rect 839 27 843 29
rect 839 21 843 23
rect 839 15 843 17
rect 839 9 843 11
rect 839 3 843 5
rect 1313 363 1317 365
rect 1313 357 1317 359
rect 1313 351 1317 353
rect 1313 345 1317 347
rect 1313 339 1317 341
rect 1313 333 1317 335
rect 1313 327 1317 329
rect 1313 321 1317 323
rect 1313 315 1317 317
rect 1313 309 1317 311
rect 1313 303 1317 305
rect 1313 297 1317 299
rect 1313 291 1317 293
rect 1313 285 1317 287
rect 1313 279 1317 281
rect 1313 273 1317 275
rect 1313 267 1317 269
rect 1313 261 1317 263
rect 1313 255 1317 257
rect 1313 249 1317 251
rect 1313 243 1317 245
rect 1313 237 1317 239
rect 1313 231 1317 233
rect 1313 225 1317 227
rect 1313 219 1317 221
rect 1313 213 1317 215
rect 1313 207 1317 209
rect 1313 201 1317 203
rect 1313 195 1317 197
rect 1313 189 1317 191
rect 1313 183 1317 185
rect 1313 177 1317 179
rect 1313 171 1317 173
rect 1313 165 1317 167
rect 1313 159 1317 161
rect 1313 153 1317 155
rect 1313 147 1317 149
rect 1313 141 1317 143
rect 1313 135 1317 137
rect 1313 129 1317 131
rect 1313 123 1317 125
rect 1313 117 1317 119
rect 1313 111 1317 113
rect 1313 105 1317 107
rect 1313 99 1317 101
rect 1313 93 1317 95
rect 1313 87 1317 89
rect 1313 81 1317 83
rect 1313 75 1317 77
rect 1313 69 1317 71
rect 1313 63 1317 65
rect 1313 57 1317 59
rect 1313 51 1317 53
rect 1313 45 1317 47
rect 1313 39 1317 41
rect 1313 33 1317 35
rect 1313 27 1317 29
rect 1313 21 1317 23
rect 1313 15 1317 17
rect 1313 9 1317 11
rect 1313 3 1317 5
rect 1787 363 1791 365
rect 1787 357 1791 359
rect 1787 351 1791 353
rect 1787 345 1791 347
rect 1787 339 1791 341
rect 1787 333 1791 335
rect 1787 327 1791 329
rect 1787 321 1791 323
rect 1787 315 1791 317
rect 1787 309 1791 311
rect 1787 303 1791 305
rect 1787 297 1791 299
rect 1787 291 1791 293
rect 1787 285 1791 287
rect 1787 279 1791 281
rect 1787 273 1791 275
rect 1787 267 1791 269
rect 1787 261 1791 263
rect 1787 255 1791 257
rect 1787 249 1791 251
rect 1787 243 1791 245
rect 1787 237 1791 239
rect 1787 231 1791 233
rect 1787 225 1791 227
rect 1787 219 1791 221
rect 1787 213 1791 215
rect 1787 207 1791 209
rect 1787 201 1791 203
rect 1787 195 1791 197
rect 1787 189 1791 191
rect 1787 183 1791 185
rect 1787 177 1791 179
rect 1787 171 1791 173
rect 1787 165 1791 167
rect 1787 159 1791 161
rect 1787 153 1791 155
rect 1787 147 1791 149
rect 1787 141 1791 143
rect 1787 135 1791 137
rect 1787 129 1791 131
rect 1787 123 1791 125
rect 1787 117 1791 119
rect 1787 111 1791 113
rect 1787 105 1791 107
rect 1787 99 1791 101
rect 1787 93 1791 95
rect 1787 87 1791 89
rect 1787 81 1791 83
rect 1787 75 1791 77
rect 1787 69 1791 71
rect 1787 63 1791 65
rect 1787 57 1791 59
rect 1787 51 1791 53
rect 1787 45 1791 47
rect 1787 39 1791 41
rect 1787 33 1791 35
rect 1787 27 1791 29
rect 1787 21 1791 23
rect 1787 15 1791 17
rect 1787 9 1791 11
rect 1787 3 1791 5
rect 2261 363 2265 365
rect 2261 357 2265 359
rect 2261 351 2265 353
rect 2261 345 2265 347
rect 2261 339 2265 341
rect 2261 333 2265 335
rect 2261 327 2265 329
rect 2261 321 2265 323
rect 2261 315 2265 317
rect 2261 309 2265 311
rect 2261 303 2265 305
rect 2261 297 2265 299
rect 2261 291 2265 293
rect 2261 285 2265 287
rect 2261 279 2265 281
rect 2261 273 2265 275
rect 2261 267 2265 269
rect 2261 261 2265 263
rect 2261 255 2265 257
rect 2261 249 2265 251
rect 2261 243 2265 245
rect 2261 237 2265 239
rect 2261 231 2265 233
rect 2261 225 2265 227
rect 2261 219 2265 221
rect 2261 213 2265 215
rect 2261 207 2265 209
rect 2261 201 2265 203
rect 2261 195 2265 197
rect 2261 189 2265 191
rect 2261 183 2265 185
rect 2261 177 2265 179
rect 2261 171 2265 173
rect 2261 165 2265 167
rect 2261 159 2265 161
rect 2261 153 2265 155
rect 2261 147 2265 149
rect 2261 141 2265 143
rect 2261 135 2265 137
rect 2261 129 2265 131
rect 2261 123 2265 125
rect 2261 117 2265 119
rect 2261 111 2265 113
rect 2261 105 2265 107
rect 2261 99 2265 101
rect 2261 93 2265 95
rect 2261 87 2265 89
rect 2261 81 2265 83
rect 2261 75 2265 77
rect 2261 69 2265 71
rect 2261 63 2265 65
rect 2261 57 2265 59
rect 2261 51 2265 53
rect 2261 45 2265 47
rect 2261 39 2265 41
rect 2261 33 2265 35
rect 2261 27 2265 29
rect 2261 21 2265 23
rect 2261 15 2265 17
rect 2261 9 2265 11
rect 2261 3 2265 5
rect 2735 363 2739 365
rect 2735 357 2739 359
rect 2735 351 2739 353
rect 2735 345 2739 347
rect 2735 339 2739 341
rect 2735 333 2739 335
rect 2735 327 2739 329
rect 2735 321 2739 323
rect 2735 315 2739 317
rect 2735 309 2739 311
rect 2735 303 2739 305
rect 2735 297 2739 299
rect 2735 291 2739 293
rect 2735 285 2739 287
rect 2735 279 2739 281
rect 2735 273 2739 275
rect 2735 267 2739 269
rect 2735 261 2739 263
rect 2735 255 2739 257
rect 2735 249 2739 251
rect 2735 243 2739 245
rect 2735 237 2739 239
rect 2735 231 2739 233
rect 2735 225 2739 227
rect 2735 219 2739 221
rect 2735 213 2739 215
rect 2735 207 2739 209
rect 2735 201 2739 203
rect 2735 195 2739 197
rect 2735 189 2739 191
rect 2735 183 2739 185
rect 2735 177 2739 179
rect 2735 171 2739 173
rect 2735 165 2739 167
rect 2735 159 2739 161
rect 2735 153 2739 155
rect 2735 147 2739 149
rect 2735 141 2739 143
rect 2735 135 2739 137
rect 2735 129 2739 131
rect 2735 123 2739 125
rect 2735 117 2739 119
rect 2735 111 2739 113
rect 2735 105 2739 107
rect 2735 99 2739 101
rect 2735 93 2739 95
rect 2735 87 2739 89
rect 2735 81 2739 83
rect 2735 75 2739 77
rect 2735 69 2739 71
rect 2735 63 2739 65
rect 2735 57 2739 59
rect 2735 51 2739 53
rect 2735 45 2739 47
rect 2735 39 2739 41
rect 2735 33 2739 35
rect 2735 27 2739 29
rect 2735 21 2739 23
rect 2735 15 2739 17
rect 2735 9 2739 11
rect 2735 3 2739 5
rect 3209 363 3213 365
rect 3209 357 3213 359
rect 3209 351 3213 353
rect 3209 345 3213 347
rect 3209 339 3213 341
rect 3209 333 3213 335
rect 3209 327 3213 329
rect 3209 321 3213 323
rect 3209 315 3213 317
rect 3209 309 3213 311
rect 3209 303 3213 305
rect 3209 297 3213 299
rect 3209 291 3213 293
rect 3209 285 3213 287
rect 3209 279 3213 281
rect 3209 273 3213 275
rect 3209 267 3213 269
rect 3209 261 3213 263
rect 3209 255 3213 257
rect 3209 249 3213 251
rect 3209 243 3213 245
rect 3209 237 3213 239
rect 3209 231 3213 233
rect 3209 225 3213 227
rect 3209 219 3213 221
rect 3209 213 3213 215
rect 3209 207 3213 209
rect 3209 201 3213 203
rect 3209 195 3213 197
rect 3209 189 3213 191
rect 3209 183 3213 185
rect 3209 177 3213 179
rect 3209 171 3213 173
rect 3209 165 3213 167
rect 3209 159 3213 161
rect 3209 153 3213 155
rect 3209 147 3213 149
rect 3209 141 3213 143
rect 3209 135 3213 137
rect 3209 129 3213 131
rect 3209 123 3213 125
rect 3209 117 3213 119
rect 3209 111 3213 113
rect 3209 105 3213 107
rect 3209 99 3213 101
rect 3209 93 3213 95
rect 3209 87 3213 89
rect 3209 81 3213 83
rect 3209 75 3213 77
rect 3209 69 3213 71
rect 3209 63 3213 65
rect 3209 57 3213 59
rect 3209 51 3213 53
rect 3209 45 3213 47
rect 3209 39 3213 41
rect 3209 33 3213 35
rect 3209 27 3213 29
rect 3209 21 3213 23
rect 3209 15 3213 17
rect 3209 9 3213 11
rect 3209 3 3213 5
rect 3683 363 3687 365
rect 3683 357 3687 359
rect 3683 351 3687 353
rect 3683 345 3687 347
rect 3683 339 3687 341
rect 3683 333 3687 335
rect 3683 327 3687 329
rect 3683 321 3687 323
rect 3683 315 3687 317
rect 3683 309 3687 311
rect 3683 303 3687 305
rect 3683 297 3687 299
rect 3683 291 3687 293
rect 3683 285 3687 287
rect 3683 279 3687 281
rect 3683 273 3687 275
rect 3683 267 3687 269
rect 3683 261 3687 263
rect 3683 255 3687 257
rect 3683 249 3687 251
rect 3683 243 3687 245
rect 3683 237 3687 239
rect 3683 231 3687 233
rect 3683 225 3687 227
rect 3683 219 3687 221
rect 3683 213 3687 215
rect 3683 207 3687 209
rect 3683 201 3687 203
rect 3683 195 3687 197
rect 3683 189 3687 191
rect 3683 183 3687 185
rect 3683 177 3687 179
rect 3683 171 3687 173
rect 3683 165 3687 167
rect 3683 159 3687 161
rect 3683 153 3687 155
rect 3683 147 3687 149
rect 3683 141 3687 143
rect 3683 135 3687 137
rect 3683 129 3687 131
rect 3683 123 3687 125
rect 3683 117 3687 119
rect 3683 111 3687 113
rect 3683 105 3687 107
rect 3683 99 3687 101
rect 3683 93 3687 95
rect 3683 87 3687 89
rect 3683 81 3687 83
rect 3683 75 3687 77
rect 3683 69 3687 71
rect 3683 63 3687 65
rect 3683 57 3687 59
rect 3683 51 3687 53
rect 3683 45 3687 47
rect 3683 39 3687 41
rect 3683 33 3687 35
rect 3683 27 3687 29
rect 3683 21 3687 23
rect 3683 15 3687 17
rect 3683 9 3687 11
rect 3683 3 3687 5
rect 4157 363 4161 365
rect 4157 357 4161 359
rect 4157 351 4161 353
rect 4157 345 4161 347
rect 4157 339 4161 341
rect 4157 333 4161 335
rect 4157 327 4161 329
rect 4157 321 4161 323
rect 4157 315 4161 317
rect 4157 309 4161 311
rect 4157 303 4161 305
rect 4157 297 4161 299
rect 4157 291 4161 293
rect 4157 285 4161 287
rect 4157 279 4161 281
rect 4157 273 4161 275
rect 4157 267 4161 269
rect 4157 261 4161 263
rect 4157 255 4161 257
rect 4157 249 4161 251
rect 4157 243 4161 245
rect 4157 237 4161 239
rect 4157 231 4161 233
rect 4157 225 4161 227
rect 4157 219 4161 221
rect 4157 213 4161 215
rect 4157 207 4161 209
rect 4157 201 4161 203
rect 4157 195 4161 197
rect 4157 189 4161 191
rect 4157 183 4161 185
rect 4157 177 4161 179
rect 4157 171 4161 173
rect 4157 165 4161 167
rect 4157 159 4161 161
rect 4157 153 4161 155
rect 4157 147 4161 149
rect 4157 141 4161 143
rect 4157 135 4161 137
rect 4157 129 4161 131
rect 4157 123 4161 125
rect 4157 117 4161 119
rect 4157 111 4161 113
rect 4157 105 4161 107
rect 4157 99 4161 101
rect 4157 93 4161 95
rect 4157 87 4161 89
rect 4157 81 4161 83
rect 4157 75 4161 77
rect 4157 69 4161 71
rect 4157 63 4161 65
rect 4157 57 4161 59
rect 4157 51 4161 53
rect 4157 45 4161 47
rect 4157 39 4161 41
rect 4157 33 4161 35
rect 4157 27 4161 29
rect 4157 21 4161 23
rect 4157 15 4161 17
rect 4157 9 4161 11
rect 4157 3 4161 5
rect 4631 363 4677 365
rect 4635 362 4677 363
rect 4635 359 4643 362
rect 4631 358 4643 359
rect 4647 358 4649 362
rect 4653 358 4655 362
rect 4659 358 4661 362
rect 4665 358 4667 362
rect 4671 358 4673 362
rect 4993 362 4997 365
rect 4631 357 4642 358
rect 4635 353 4638 357
rect 4631 351 4642 353
rect 4635 347 4638 351
rect 4631 345 4642 347
rect 4635 341 4638 345
rect 4631 339 4642 341
rect 4635 335 4638 339
rect 4631 333 4642 335
rect 4635 329 4638 333
rect 4631 327 4642 329
rect 4635 323 4638 327
rect 4993 356 4997 358
rect 4993 350 4997 352
rect 4993 344 4997 346
rect 4993 338 4997 340
rect 4993 332 4997 334
rect 4993 326 4997 328
rect 4631 321 4635 323
rect 4631 315 4635 317
rect 4993 320 4997 322
rect 4631 309 4635 311
rect 4631 303 4635 305
rect 4631 297 4635 299
rect 4631 291 4635 293
rect 4631 285 4635 287
rect 4631 279 4635 281
rect 4631 273 4635 275
rect 4631 267 4635 269
rect 4631 261 4635 263
rect 4631 255 4635 257
rect 4631 249 4635 251
rect 4631 243 4635 245
rect 4631 237 4635 239
rect 4631 231 4635 233
rect 4631 225 4635 227
rect 4631 219 4635 221
rect 4644 259 4680 260
rect 4644 255 4645 259
rect 4649 255 4657 259
rect 4661 255 4669 259
rect 4673 255 4680 259
rect 4644 253 4680 255
rect 4644 249 4645 253
rect 4649 249 4651 253
rect 4655 249 4657 253
rect 4661 249 4663 253
rect 4667 249 4669 253
rect 4673 249 4675 253
rect 4679 249 4680 253
rect 4644 247 4680 249
rect 4644 243 4651 247
rect 4655 243 4663 247
rect 4667 243 4675 247
rect 4679 243 4680 247
rect 4644 241 4680 243
rect 4644 237 4645 241
rect 4649 237 4651 241
rect 4655 237 4657 241
rect 4661 237 4663 241
rect 4667 237 4669 241
rect 4673 237 4675 241
rect 4679 237 4680 241
rect 4644 235 4680 237
rect 4644 231 4645 235
rect 4649 231 4657 235
rect 4661 231 4669 235
rect 4673 231 4680 235
rect 4644 229 4680 231
rect 4644 225 4645 229
rect 4649 225 4651 229
rect 4655 225 4657 229
rect 4661 225 4663 229
rect 4667 225 4669 229
rect 4673 225 4675 229
rect 4679 225 4680 229
rect 4644 223 4680 225
rect 4644 219 4651 223
rect 4655 219 4663 223
rect 4667 219 4675 223
rect 4679 219 4680 223
rect 4644 218 4680 219
rect 4631 213 4635 215
rect 4631 207 4635 209
rect 4631 201 4635 203
rect 4631 195 4635 197
rect 4631 189 4635 191
rect 4631 183 4635 185
rect 4631 177 4635 179
rect 4631 171 4635 173
rect 4631 165 4635 167
rect 4631 159 4635 161
rect 4631 153 4635 155
rect 4631 147 4635 149
rect 4631 141 4635 143
rect 4631 135 4635 137
rect 4631 129 4635 131
rect 4631 123 4635 125
rect 4631 117 4635 119
rect 4631 111 4635 113
rect 4631 105 4635 107
rect 4631 99 4635 101
rect 4631 93 4635 95
rect 4631 87 4635 89
rect 4631 81 4635 83
rect 4631 75 4635 77
rect 4631 69 4635 71
rect 4631 63 4635 65
rect 4631 57 4635 59
rect 4631 51 4635 53
rect 4631 45 4635 47
rect 4631 39 4635 41
rect 4631 33 4635 35
rect 4631 27 4635 29
rect 4631 21 4635 23
rect 4631 15 4635 17
rect 4631 9 4635 11
rect 4635 5 4638 7
rect 4631 3 4638 5
rect 4642 3 4644 7
rect 4648 3 4650 7
rect 4654 3 4656 7
rect 4660 3 4662 7
rect 4666 3 4668 7
rect 4672 3 4674 7
rect 4678 3 4680 7
<< m2contact >>
rect 539 509 543 513
rect 545 509 549 513
rect 551 509 555 513
rect 557 509 561 513
rect 563 509 567 513
rect 569 509 573 513
rect 575 509 579 513
rect 539 495 543 499
rect 545 495 549 499
rect 551 495 555 499
rect 557 495 561 499
rect 563 495 567 499
rect 569 495 573 499
rect 575 495 579 499
rect 539 483 543 487
rect 545 483 549 487
rect 551 483 555 487
rect 557 483 561 487
rect 563 483 567 487
rect 569 483 573 487
rect 575 483 579 487
rect 539 477 543 481
rect 545 477 549 481
rect 551 477 555 481
rect 557 477 561 481
rect 563 477 567 481
rect 569 477 573 481
rect 575 477 579 481
rect 539 466 543 470
rect 545 466 549 470
rect 551 466 555 470
rect 557 466 561 470
rect 563 466 567 470
rect 569 466 573 470
rect 575 466 579 470
rect 583 509 592 513
rect 495 441 499 450
rect 501 441 505 450
rect 507 441 511 450
rect 513 441 517 450
rect 519 441 523 450
rect 525 441 529 450
rect 531 441 535 450
rect 495 435 499 439
rect 501 435 505 439
rect 507 435 511 439
rect 513 435 517 439
rect 519 435 523 439
rect 525 435 529 439
rect 531 435 535 439
rect 495 429 499 433
rect 501 429 505 433
rect 507 429 511 433
rect 513 429 517 433
rect 519 429 523 433
rect 525 429 529 433
rect 531 429 535 433
rect 495 423 499 427
rect 501 423 505 427
rect 507 423 511 427
rect 513 423 517 427
rect 519 423 523 427
rect 525 423 529 427
rect 531 423 535 427
rect 495 412 499 421
rect 501 412 505 421
rect 507 412 511 421
rect 513 412 517 421
rect 519 412 523 421
rect 525 412 529 421
rect 531 412 535 421
rect 578 456 582 460
rect 588 456 592 460
rect 616 509 625 513
rect 629 509 633 513
rect 635 509 639 513
rect 641 509 645 513
rect 647 509 651 513
rect 653 509 657 513
rect 659 509 663 513
rect 665 509 669 513
rect 629 495 633 499
rect 635 495 639 499
rect 641 495 645 499
rect 647 495 651 499
rect 653 495 657 499
rect 659 495 663 499
rect 629 483 633 487
rect 635 483 639 487
rect 641 483 645 487
rect 647 483 651 487
rect 653 483 657 487
rect 659 483 663 487
rect 665 483 669 487
rect 629 477 633 481
rect 635 477 639 481
rect 641 477 645 481
rect 647 477 651 481
rect 653 477 657 481
rect 659 477 663 481
rect 665 477 669 481
rect 629 466 633 470
rect 635 466 639 470
rect 641 466 645 470
rect 647 466 651 470
rect 653 466 657 470
rect 659 466 663 470
rect 665 466 669 470
rect 616 456 620 460
rect 626 456 630 460
rect 673 509 677 513
rect 679 509 683 513
rect 685 509 689 513
rect 691 509 695 513
rect 697 509 701 513
rect 703 509 707 513
rect 709 509 713 513
rect 673 441 677 450
rect 679 441 683 450
rect 685 441 689 450
rect 691 441 695 450
rect 697 441 701 450
rect 703 441 707 450
rect 709 441 713 450
rect 673 435 677 439
rect 679 435 683 439
rect 685 435 689 439
rect 691 435 695 439
rect 697 435 701 439
rect 703 435 707 439
rect 709 435 713 439
rect 673 429 677 433
rect 679 429 683 433
rect 685 429 689 433
rect 691 429 695 433
rect 697 429 701 433
rect 703 429 707 433
rect 709 429 713 433
rect 673 423 677 427
rect 679 423 683 427
rect 685 423 689 427
rect 691 423 695 427
rect 697 423 701 427
rect 703 423 707 427
rect 709 423 713 427
rect 673 412 677 421
rect 679 412 683 421
rect 685 412 689 421
rect 691 412 695 421
rect 697 412 701 421
rect 703 412 707 421
rect 709 412 713 421
rect 539 402 543 406
rect 545 402 549 406
rect 551 402 555 406
rect 557 402 561 406
rect 563 402 567 406
rect 569 402 573 406
rect 575 402 579 406
rect 539 390 543 394
rect 545 390 549 394
rect 551 390 555 394
rect 557 390 561 394
rect 563 390 567 394
rect 569 390 573 394
rect 575 390 579 394
rect 545 378 549 382
rect 551 378 555 382
rect 557 378 561 382
rect 563 378 567 382
rect 569 378 573 382
rect 575 378 579 382
rect 629 402 633 406
rect 635 402 639 406
rect 641 402 645 406
rect 647 402 651 406
rect 653 402 657 406
rect 659 402 663 406
rect 665 402 669 406
rect 629 390 633 394
rect 635 390 639 394
rect 641 390 645 394
rect 647 390 651 394
rect 653 390 657 394
rect 659 390 663 394
rect 665 390 669 394
rect 629 378 633 382
rect 635 378 639 382
rect 641 378 645 382
rect 647 378 651 382
rect 653 378 657 382
rect 659 378 663 382
rect 969 509 973 513
rect 975 509 979 513
rect 981 509 985 513
rect 987 509 991 513
rect 993 509 997 513
rect 999 509 1003 513
rect 1005 509 1009 513
rect 969 441 973 450
rect 975 441 979 450
rect 981 441 985 450
rect 987 441 991 450
rect 993 441 997 450
rect 999 441 1003 450
rect 1005 441 1009 450
rect 969 435 973 439
rect 975 435 979 439
rect 981 435 985 439
rect 987 435 991 439
rect 993 435 997 439
rect 999 435 1003 439
rect 1005 435 1009 439
rect 969 429 973 433
rect 975 429 979 433
rect 981 429 985 433
rect 987 429 991 433
rect 993 429 997 433
rect 999 429 1003 433
rect 1005 429 1009 433
rect 969 423 973 427
rect 975 423 979 427
rect 981 423 985 427
rect 987 423 991 427
rect 993 423 997 427
rect 999 423 1003 427
rect 1005 423 1009 427
rect 969 412 973 421
rect 975 412 979 421
rect 981 412 985 421
rect 987 412 991 421
rect 993 412 997 421
rect 999 412 1003 421
rect 1005 412 1009 421
rect 1013 509 1017 513
rect 1019 509 1023 513
rect 1025 509 1029 513
rect 1031 509 1035 513
rect 1037 509 1041 513
rect 1043 509 1047 513
rect 1049 509 1053 513
rect 1019 495 1023 499
rect 1025 495 1029 499
rect 1031 495 1035 499
rect 1037 495 1041 499
rect 1043 495 1047 499
rect 1049 495 1053 499
rect 1013 483 1017 487
rect 1019 483 1023 487
rect 1025 483 1029 487
rect 1031 483 1035 487
rect 1037 483 1041 487
rect 1043 483 1047 487
rect 1049 483 1053 487
rect 1013 477 1017 481
rect 1019 477 1023 481
rect 1025 477 1029 481
rect 1031 477 1035 481
rect 1037 477 1041 481
rect 1043 477 1047 481
rect 1049 477 1053 481
rect 1013 465 1017 469
rect 1019 465 1023 469
rect 1025 465 1029 469
rect 1031 465 1035 469
rect 1037 465 1041 469
rect 1043 465 1047 469
rect 1049 465 1053 469
rect 1057 509 1066 513
rect 1052 456 1056 460
rect 1062 456 1066 460
rect 1090 509 1099 513
rect 1103 509 1107 513
rect 1109 509 1113 513
rect 1115 509 1119 513
rect 1121 509 1125 513
rect 1127 509 1131 513
rect 1133 509 1137 513
rect 1139 509 1143 513
rect 1103 495 1107 499
rect 1109 495 1113 499
rect 1115 495 1119 499
rect 1121 495 1125 499
rect 1127 495 1131 499
rect 1133 495 1137 499
rect 1103 483 1107 487
rect 1109 483 1113 487
rect 1115 483 1119 487
rect 1121 483 1125 487
rect 1127 483 1131 487
rect 1133 483 1137 487
rect 1139 483 1143 487
rect 1103 477 1107 481
rect 1109 477 1113 481
rect 1115 477 1119 481
rect 1121 477 1125 481
rect 1127 477 1131 481
rect 1133 477 1137 481
rect 1139 477 1143 481
rect 1103 465 1107 469
rect 1109 465 1113 469
rect 1115 465 1119 469
rect 1121 465 1125 469
rect 1127 465 1131 469
rect 1133 465 1137 469
rect 1139 465 1143 469
rect 1090 456 1094 460
rect 1100 456 1104 460
rect 1147 509 1151 513
rect 1153 509 1157 513
rect 1159 509 1163 513
rect 1165 509 1169 513
rect 1171 509 1175 513
rect 1177 509 1181 513
rect 1183 509 1187 513
rect 1147 441 1151 450
rect 1153 441 1157 450
rect 1159 441 1163 450
rect 1165 441 1169 450
rect 1171 441 1175 450
rect 1177 441 1181 450
rect 1183 441 1187 450
rect 1147 435 1151 439
rect 1153 435 1157 439
rect 1159 435 1163 439
rect 1165 435 1169 439
rect 1171 435 1175 439
rect 1177 435 1181 439
rect 1183 435 1187 439
rect 1147 429 1151 433
rect 1153 429 1157 433
rect 1159 429 1163 433
rect 1165 429 1169 433
rect 1171 429 1175 433
rect 1177 429 1181 433
rect 1183 429 1187 433
rect 1147 423 1151 427
rect 1153 423 1157 427
rect 1159 423 1163 427
rect 1165 423 1169 427
rect 1171 423 1175 427
rect 1177 423 1181 427
rect 1183 423 1187 427
rect 1147 412 1151 421
rect 1153 412 1157 421
rect 1159 412 1163 421
rect 1165 412 1169 421
rect 1171 412 1175 421
rect 1177 412 1181 421
rect 1183 412 1187 421
rect 1013 402 1017 406
rect 1019 402 1023 406
rect 1025 402 1029 406
rect 1031 402 1035 406
rect 1037 402 1041 406
rect 1043 402 1047 406
rect 1049 402 1053 406
rect 1013 390 1017 394
rect 1019 390 1023 394
rect 1025 390 1029 394
rect 1031 390 1035 394
rect 1037 390 1041 394
rect 1043 390 1047 394
rect 1049 390 1053 394
rect 1019 378 1023 382
rect 1025 378 1029 382
rect 1031 378 1035 382
rect 1037 378 1041 382
rect 1043 378 1047 382
rect 1049 378 1053 382
rect 1103 402 1107 406
rect 1109 402 1113 406
rect 1115 402 1119 406
rect 1121 402 1125 406
rect 1127 402 1131 406
rect 1133 402 1137 406
rect 1139 402 1143 406
rect 1103 390 1107 394
rect 1109 390 1113 394
rect 1115 390 1119 394
rect 1121 390 1125 394
rect 1127 390 1131 394
rect 1133 390 1137 394
rect 1139 390 1143 394
rect 1103 378 1107 382
rect 1109 378 1113 382
rect 1115 378 1119 382
rect 1121 378 1125 382
rect 1127 378 1131 382
rect 1133 378 1137 382
rect 1443 509 1447 513
rect 1449 509 1453 513
rect 1455 509 1459 513
rect 1461 509 1465 513
rect 1467 509 1471 513
rect 1473 509 1477 513
rect 1479 509 1483 513
rect 1443 441 1447 450
rect 1449 441 1453 450
rect 1455 441 1459 450
rect 1461 441 1465 450
rect 1467 441 1471 450
rect 1473 441 1477 450
rect 1479 441 1483 450
rect 1443 435 1447 439
rect 1449 435 1453 439
rect 1455 435 1459 439
rect 1461 435 1465 439
rect 1467 435 1471 439
rect 1473 435 1477 439
rect 1479 435 1483 439
rect 1443 429 1447 433
rect 1449 429 1453 433
rect 1455 429 1459 433
rect 1461 429 1465 433
rect 1467 429 1471 433
rect 1473 429 1477 433
rect 1479 429 1483 433
rect 1443 423 1447 427
rect 1449 423 1453 427
rect 1455 423 1459 427
rect 1461 423 1465 427
rect 1467 423 1471 427
rect 1473 423 1477 427
rect 1479 423 1483 427
rect 1443 412 1447 421
rect 1449 412 1453 421
rect 1455 412 1459 421
rect 1461 412 1465 421
rect 1467 412 1471 421
rect 1473 412 1477 421
rect 1479 412 1483 421
rect 1487 509 1491 513
rect 1493 509 1497 513
rect 1499 509 1503 513
rect 1505 509 1509 513
rect 1511 509 1515 513
rect 1517 509 1521 513
rect 1523 509 1527 513
rect 1493 495 1497 499
rect 1499 495 1503 499
rect 1505 495 1509 499
rect 1511 495 1515 499
rect 1517 495 1521 499
rect 1523 495 1527 499
rect 1487 483 1491 487
rect 1493 483 1497 487
rect 1499 483 1503 487
rect 1505 483 1509 487
rect 1511 483 1515 487
rect 1517 483 1521 487
rect 1523 483 1527 487
rect 1487 477 1491 481
rect 1493 477 1497 481
rect 1499 477 1503 481
rect 1505 477 1509 481
rect 1511 477 1515 481
rect 1517 477 1521 481
rect 1523 477 1527 481
rect 1487 465 1491 469
rect 1493 465 1497 469
rect 1499 465 1503 469
rect 1505 465 1509 469
rect 1511 465 1515 469
rect 1517 465 1521 469
rect 1523 465 1527 469
rect 1531 509 1540 513
rect 1526 456 1530 460
rect 1536 456 1540 460
rect 1564 509 1573 513
rect 1577 509 1581 513
rect 1583 509 1587 513
rect 1589 509 1593 513
rect 1595 509 1599 513
rect 1601 509 1605 513
rect 1607 509 1611 513
rect 1613 509 1617 513
rect 1577 495 1581 499
rect 1583 495 1587 499
rect 1589 495 1593 499
rect 1595 495 1599 499
rect 1601 495 1605 499
rect 1607 495 1611 499
rect 1577 483 1581 487
rect 1583 483 1587 487
rect 1589 483 1593 487
rect 1595 483 1599 487
rect 1601 483 1605 487
rect 1607 483 1611 487
rect 1613 483 1617 487
rect 1577 477 1581 481
rect 1583 477 1587 481
rect 1589 477 1593 481
rect 1595 477 1599 481
rect 1601 477 1605 481
rect 1607 477 1611 481
rect 1613 477 1617 481
rect 1577 465 1581 469
rect 1583 465 1587 469
rect 1589 465 1593 469
rect 1595 465 1599 469
rect 1601 465 1605 469
rect 1607 465 1611 469
rect 1613 465 1617 469
rect 1564 456 1568 460
rect 1574 456 1578 460
rect 1621 509 1625 513
rect 1627 509 1631 513
rect 1633 509 1637 513
rect 1639 509 1643 513
rect 1645 509 1649 513
rect 1651 509 1655 513
rect 1657 509 1661 513
rect 1621 441 1625 450
rect 1627 441 1631 450
rect 1633 441 1637 450
rect 1639 441 1643 450
rect 1645 441 1649 450
rect 1651 441 1655 450
rect 1657 441 1661 450
rect 1621 435 1625 439
rect 1627 435 1631 439
rect 1633 435 1637 439
rect 1639 435 1643 439
rect 1645 435 1649 439
rect 1651 435 1655 439
rect 1657 435 1661 439
rect 1621 429 1625 433
rect 1627 429 1631 433
rect 1633 429 1637 433
rect 1639 429 1643 433
rect 1645 429 1649 433
rect 1651 429 1655 433
rect 1657 429 1661 433
rect 1621 423 1625 427
rect 1627 423 1631 427
rect 1633 423 1637 427
rect 1639 423 1643 427
rect 1645 423 1649 427
rect 1651 423 1655 427
rect 1657 423 1661 427
rect 1621 412 1625 421
rect 1627 412 1631 421
rect 1633 412 1637 421
rect 1639 412 1643 421
rect 1645 412 1649 421
rect 1651 412 1655 421
rect 1657 412 1661 421
rect 1487 402 1491 406
rect 1493 402 1497 406
rect 1499 402 1503 406
rect 1505 402 1509 406
rect 1511 402 1515 406
rect 1517 402 1521 406
rect 1523 402 1527 406
rect 1487 390 1491 394
rect 1493 390 1497 394
rect 1499 390 1503 394
rect 1505 390 1509 394
rect 1511 390 1515 394
rect 1517 390 1521 394
rect 1523 390 1527 394
rect 1493 378 1497 382
rect 1499 378 1503 382
rect 1505 378 1509 382
rect 1511 378 1515 382
rect 1517 378 1521 382
rect 1523 378 1527 382
rect 1577 402 1581 406
rect 1583 402 1587 406
rect 1589 402 1593 406
rect 1595 402 1599 406
rect 1601 402 1605 406
rect 1607 402 1611 406
rect 1613 402 1617 406
rect 1577 390 1581 394
rect 1583 390 1587 394
rect 1589 390 1593 394
rect 1595 390 1599 394
rect 1601 390 1605 394
rect 1607 390 1611 394
rect 1613 390 1617 394
rect 1577 378 1581 382
rect 1583 378 1587 382
rect 1589 378 1593 382
rect 1595 378 1599 382
rect 1601 378 1605 382
rect 1607 378 1611 382
rect 1917 509 1921 513
rect 1923 509 1927 513
rect 1929 509 1933 513
rect 1935 509 1939 513
rect 1941 509 1945 513
rect 1947 509 1951 513
rect 1953 509 1957 513
rect 1917 441 1921 450
rect 1923 441 1927 450
rect 1929 441 1933 450
rect 1935 441 1939 450
rect 1941 441 1945 450
rect 1947 441 1951 450
rect 1953 441 1957 450
rect 1917 435 1921 439
rect 1923 435 1927 439
rect 1929 435 1933 439
rect 1935 435 1939 439
rect 1941 435 1945 439
rect 1947 435 1951 439
rect 1953 435 1957 439
rect 1917 429 1921 433
rect 1923 429 1927 433
rect 1929 429 1933 433
rect 1935 429 1939 433
rect 1941 429 1945 433
rect 1947 429 1951 433
rect 1953 429 1957 433
rect 1917 423 1921 427
rect 1923 423 1927 427
rect 1929 423 1933 427
rect 1935 423 1939 427
rect 1941 423 1945 427
rect 1947 423 1951 427
rect 1953 423 1957 427
rect 1917 412 1921 421
rect 1923 412 1927 421
rect 1929 412 1933 421
rect 1935 412 1939 421
rect 1941 412 1945 421
rect 1947 412 1951 421
rect 1953 412 1957 421
rect 1961 509 1965 513
rect 1967 509 1971 513
rect 1973 509 1977 513
rect 1979 509 1983 513
rect 1985 509 1989 513
rect 1991 509 1995 513
rect 1997 509 2001 513
rect 1967 495 1971 499
rect 1973 495 1977 499
rect 1979 495 1983 499
rect 1985 495 1989 499
rect 1991 495 1995 499
rect 1997 495 2001 499
rect 1961 483 1965 487
rect 1967 483 1971 487
rect 1973 483 1977 487
rect 1979 483 1983 487
rect 1985 483 1989 487
rect 1991 483 1995 487
rect 1997 483 2001 487
rect 1961 477 1965 481
rect 1967 477 1971 481
rect 1973 477 1977 481
rect 1979 477 1983 481
rect 1985 477 1989 481
rect 1991 477 1995 481
rect 1997 477 2001 481
rect 1961 465 1965 469
rect 1967 465 1971 469
rect 1973 465 1977 469
rect 1979 465 1983 469
rect 1985 465 1989 469
rect 1991 465 1995 469
rect 1997 465 2001 469
rect 2005 509 2014 513
rect 2000 456 2004 460
rect 2010 456 2014 460
rect 2038 509 2047 513
rect 2051 509 2055 513
rect 2057 509 2061 513
rect 2063 509 2067 513
rect 2069 509 2073 513
rect 2075 509 2079 513
rect 2081 509 2085 513
rect 2087 509 2091 513
rect 2051 495 2055 499
rect 2057 495 2061 499
rect 2063 495 2067 499
rect 2069 495 2073 499
rect 2075 495 2079 499
rect 2081 495 2085 499
rect 2051 483 2055 487
rect 2057 483 2061 487
rect 2063 483 2067 487
rect 2069 483 2073 487
rect 2075 483 2079 487
rect 2081 483 2085 487
rect 2087 483 2091 487
rect 2051 477 2055 481
rect 2057 477 2061 481
rect 2063 477 2067 481
rect 2069 477 2073 481
rect 2075 477 2079 481
rect 2081 477 2085 481
rect 2087 477 2091 481
rect 2051 465 2055 469
rect 2057 465 2061 469
rect 2063 465 2067 469
rect 2069 465 2073 469
rect 2075 465 2079 469
rect 2081 465 2085 469
rect 2087 465 2091 469
rect 2038 456 2042 460
rect 2048 456 2052 460
rect 2095 509 2099 513
rect 2101 509 2105 513
rect 2107 509 2111 513
rect 2113 509 2117 513
rect 2119 509 2123 513
rect 2125 509 2129 513
rect 2131 509 2135 513
rect 2095 441 2099 450
rect 2101 441 2105 450
rect 2107 441 2111 450
rect 2113 441 2117 450
rect 2119 441 2123 450
rect 2125 441 2129 450
rect 2131 441 2135 450
rect 2095 435 2099 439
rect 2101 435 2105 439
rect 2107 435 2111 439
rect 2113 435 2117 439
rect 2119 435 2123 439
rect 2125 435 2129 439
rect 2131 435 2135 439
rect 2095 429 2099 433
rect 2101 429 2105 433
rect 2107 429 2111 433
rect 2113 429 2117 433
rect 2119 429 2123 433
rect 2125 429 2129 433
rect 2131 429 2135 433
rect 2095 423 2099 427
rect 2101 423 2105 427
rect 2107 423 2111 427
rect 2113 423 2117 427
rect 2119 423 2123 427
rect 2125 423 2129 427
rect 2131 423 2135 427
rect 2095 412 2099 421
rect 2101 412 2105 421
rect 2107 412 2111 421
rect 2113 412 2117 421
rect 2119 412 2123 421
rect 2125 412 2129 421
rect 2131 412 2135 421
rect 1961 402 1965 406
rect 1967 402 1971 406
rect 1973 402 1977 406
rect 1979 402 1983 406
rect 1985 402 1989 406
rect 1991 402 1995 406
rect 1997 402 2001 406
rect 1961 390 1965 394
rect 1967 390 1971 394
rect 1973 390 1977 394
rect 1979 390 1983 394
rect 1985 390 1989 394
rect 1991 390 1995 394
rect 1997 390 2001 394
rect 1967 378 1971 382
rect 1973 378 1977 382
rect 1979 378 1983 382
rect 1985 378 1989 382
rect 1991 378 1995 382
rect 1997 378 2001 382
rect 2051 402 2055 406
rect 2057 402 2061 406
rect 2063 402 2067 406
rect 2069 402 2073 406
rect 2075 402 2079 406
rect 2081 402 2085 406
rect 2087 402 2091 406
rect 2051 390 2055 394
rect 2057 390 2061 394
rect 2063 390 2067 394
rect 2069 390 2073 394
rect 2075 390 2079 394
rect 2081 390 2085 394
rect 2087 390 2091 394
rect 2051 378 2055 382
rect 2057 378 2061 382
rect 2063 378 2067 382
rect 2069 378 2073 382
rect 2075 378 2079 382
rect 2081 378 2085 382
rect 2391 509 2395 513
rect 2397 509 2401 513
rect 2403 509 2407 513
rect 2409 509 2413 513
rect 2415 509 2419 513
rect 2421 509 2425 513
rect 2427 509 2431 513
rect 2391 441 2395 450
rect 2397 441 2401 450
rect 2403 441 2407 450
rect 2409 441 2413 450
rect 2415 441 2419 450
rect 2421 441 2425 450
rect 2427 441 2431 450
rect 2391 435 2395 439
rect 2397 435 2401 439
rect 2403 435 2407 439
rect 2409 435 2413 439
rect 2415 435 2419 439
rect 2421 435 2425 439
rect 2427 435 2431 439
rect 2391 429 2395 433
rect 2397 429 2401 433
rect 2403 429 2407 433
rect 2409 429 2413 433
rect 2415 429 2419 433
rect 2421 429 2425 433
rect 2427 429 2431 433
rect 2391 423 2395 427
rect 2397 423 2401 427
rect 2403 423 2407 427
rect 2409 423 2413 427
rect 2415 423 2419 427
rect 2421 423 2425 427
rect 2427 423 2431 427
rect 2391 412 2395 421
rect 2397 412 2401 421
rect 2403 412 2407 421
rect 2409 412 2413 421
rect 2415 412 2419 421
rect 2421 412 2425 421
rect 2427 412 2431 421
rect 2435 509 2439 513
rect 2441 509 2445 513
rect 2447 509 2451 513
rect 2453 509 2457 513
rect 2459 509 2463 513
rect 2465 509 2469 513
rect 2471 509 2475 513
rect 2441 495 2445 499
rect 2447 495 2451 499
rect 2453 495 2457 499
rect 2459 495 2463 499
rect 2465 495 2469 499
rect 2471 495 2475 499
rect 2435 483 2439 487
rect 2441 483 2445 487
rect 2447 483 2451 487
rect 2453 483 2457 487
rect 2459 483 2463 487
rect 2465 483 2469 487
rect 2471 483 2475 487
rect 2435 477 2439 481
rect 2441 477 2445 481
rect 2447 477 2451 481
rect 2453 477 2457 481
rect 2459 477 2463 481
rect 2465 477 2469 481
rect 2471 477 2475 481
rect 2435 465 2439 469
rect 2441 465 2445 469
rect 2447 465 2451 469
rect 2453 465 2457 469
rect 2459 465 2463 469
rect 2465 465 2469 469
rect 2471 465 2475 469
rect 2479 509 2488 513
rect 2474 456 2478 460
rect 2484 456 2488 460
rect 2512 509 2521 513
rect 2525 509 2529 513
rect 2531 509 2535 513
rect 2537 509 2541 513
rect 2543 509 2547 513
rect 2549 509 2553 513
rect 2555 509 2559 513
rect 2561 509 2565 513
rect 2525 495 2529 499
rect 2531 495 2535 499
rect 2537 495 2541 499
rect 2543 495 2547 499
rect 2549 495 2553 499
rect 2555 495 2559 499
rect 2525 483 2529 487
rect 2531 483 2535 487
rect 2537 483 2541 487
rect 2543 483 2547 487
rect 2549 483 2553 487
rect 2555 483 2559 487
rect 2561 483 2565 487
rect 2525 477 2529 481
rect 2531 477 2535 481
rect 2537 477 2541 481
rect 2543 477 2547 481
rect 2549 477 2553 481
rect 2555 477 2559 481
rect 2561 477 2565 481
rect 2525 465 2529 469
rect 2531 465 2535 469
rect 2537 465 2541 469
rect 2543 465 2547 469
rect 2549 465 2553 469
rect 2555 465 2559 469
rect 2561 465 2565 469
rect 2512 456 2516 460
rect 2522 456 2526 460
rect 2569 509 2573 513
rect 2575 509 2579 513
rect 2581 509 2585 513
rect 2587 509 2591 513
rect 2593 509 2597 513
rect 2599 509 2603 513
rect 2605 509 2609 513
rect 2569 441 2573 450
rect 2575 441 2579 450
rect 2581 441 2585 450
rect 2587 441 2591 450
rect 2593 441 2597 450
rect 2599 441 2603 450
rect 2605 441 2609 450
rect 2569 435 2573 439
rect 2575 435 2579 439
rect 2581 435 2585 439
rect 2587 435 2591 439
rect 2593 435 2597 439
rect 2599 435 2603 439
rect 2605 435 2609 439
rect 2569 429 2573 433
rect 2575 429 2579 433
rect 2581 429 2585 433
rect 2587 429 2591 433
rect 2593 429 2597 433
rect 2599 429 2603 433
rect 2605 429 2609 433
rect 2569 423 2573 427
rect 2575 423 2579 427
rect 2581 423 2585 427
rect 2587 423 2591 427
rect 2593 423 2597 427
rect 2599 423 2603 427
rect 2605 423 2609 427
rect 2569 412 2573 421
rect 2575 412 2579 421
rect 2581 412 2585 421
rect 2587 412 2591 421
rect 2593 412 2597 421
rect 2599 412 2603 421
rect 2605 412 2609 421
rect 2435 402 2439 406
rect 2441 402 2445 406
rect 2447 402 2451 406
rect 2453 402 2457 406
rect 2459 402 2463 406
rect 2465 402 2469 406
rect 2471 402 2475 406
rect 2435 390 2439 394
rect 2441 390 2445 394
rect 2447 390 2451 394
rect 2453 390 2457 394
rect 2459 390 2463 394
rect 2465 390 2469 394
rect 2471 390 2475 394
rect 2441 378 2445 382
rect 2447 378 2451 382
rect 2453 378 2457 382
rect 2459 378 2463 382
rect 2465 378 2469 382
rect 2471 378 2475 382
rect 2525 402 2529 406
rect 2531 402 2535 406
rect 2537 402 2541 406
rect 2543 402 2547 406
rect 2549 402 2553 406
rect 2555 402 2559 406
rect 2561 402 2565 406
rect 2525 390 2529 394
rect 2531 390 2535 394
rect 2537 390 2541 394
rect 2543 390 2547 394
rect 2549 390 2553 394
rect 2555 390 2559 394
rect 2561 390 2565 394
rect 2525 378 2529 382
rect 2531 378 2535 382
rect 2537 378 2541 382
rect 2543 378 2547 382
rect 2549 378 2553 382
rect 2555 378 2559 382
rect 2865 509 2869 513
rect 2871 509 2875 513
rect 2877 509 2881 513
rect 2883 509 2887 513
rect 2889 509 2893 513
rect 2895 509 2899 513
rect 2901 509 2905 513
rect 2865 441 2869 450
rect 2871 441 2875 450
rect 2877 441 2881 450
rect 2883 441 2887 450
rect 2889 441 2893 450
rect 2895 441 2899 450
rect 2901 441 2905 450
rect 2865 435 2869 439
rect 2871 435 2875 439
rect 2877 435 2881 439
rect 2883 435 2887 439
rect 2889 435 2893 439
rect 2895 435 2899 439
rect 2901 435 2905 439
rect 2865 429 2869 433
rect 2871 429 2875 433
rect 2877 429 2881 433
rect 2883 429 2887 433
rect 2889 429 2893 433
rect 2895 429 2899 433
rect 2901 429 2905 433
rect 2865 423 2869 427
rect 2871 423 2875 427
rect 2877 423 2881 427
rect 2883 423 2887 427
rect 2889 423 2893 427
rect 2895 423 2899 427
rect 2901 423 2905 427
rect 2865 412 2869 421
rect 2871 412 2875 421
rect 2877 412 2881 421
rect 2883 412 2887 421
rect 2889 412 2893 421
rect 2895 412 2899 421
rect 2901 412 2905 421
rect 2909 509 2913 513
rect 2915 509 2919 513
rect 2921 509 2925 513
rect 2927 509 2931 513
rect 2933 509 2937 513
rect 2939 509 2943 513
rect 2945 509 2949 513
rect 2915 495 2919 499
rect 2921 495 2925 499
rect 2927 495 2931 499
rect 2933 495 2937 499
rect 2939 495 2943 499
rect 2945 495 2949 499
rect 2909 483 2913 487
rect 2915 483 2919 487
rect 2921 483 2925 487
rect 2927 483 2931 487
rect 2933 483 2937 487
rect 2939 483 2943 487
rect 2945 483 2949 487
rect 2909 477 2913 481
rect 2915 477 2919 481
rect 2921 477 2925 481
rect 2927 477 2931 481
rect 2933 477 2937 481
rect 2939 477 2943 481
rect 2945 477 2949 481
rect 2909 465 2913 469
rect 2915 465 2919 469
rect 2921 465 2925 469
rect 2927 465 2931 469
rect 2933 465 2937 469
rect 2939 465 2943 469
rect 2945 465 2949 469
rect 2953 509 2962 513
rect 2948 456 2952 460
rect 2958 456 2962 460
rect 2986 509 2995 513
rect 2999 509 3003 513
rect 3005 509 3009 513
rect 3011 509 3015 513
rect 3017 509 3021 513
rect 3023 509 3027 513
rect 3029 509 3033 513
rect 3035 509 3039 513
rect 2999 495 3003 499
rect 3005 495 3009 499
rect 3011 495 3015 499
rect 3017 495 3021 499
rect 3023 495 3027 499
rect 3029 495 3033 499
rect 2999 483 3003 487
rect 3005 483 3009 487
rect 3011 483 3015 487
rect 3017 483 3021 487
rect 3023 483 3027 487
rect 3029 483 3033 487
rect 3035 483 3039 487
rect 2999 477 3003 481
rect 3005 477 3009 481
rect 3011 477 3015 481
rect 3017 477 3021 481
rect 3023 477 3027 481
rect 3029 477 3033 481
rect 3035 477 3039 481
rect 2999 465 3003 469
rect 3005 465 3009 469
rect 3011 465 3015 469
rect 3017 465 3021 469
rect 3023 465 3027 469
rect 3029 465 3033 469
rect 3035 465 3039 469
rect 2986 456 2990 460
rect 2996 456 3000 460
rect 3043 509 3047 513
rect 3049 509 3053 513
rect 3055 509 3059 513
rect 3061 509 3065 513
rect 3067 509 3071 513
rect 3073 509 3077 513
rect 3079 509 3083 513
rect 3043 441 3047 450
rect 3049 441 3053 450
rect 3055 441 3059 450
rect 3061 441 3065 450
rect 3067 441 3071 450
rect 3073 441 3077 450
rect 3079 441 3083 450
rect 3043 435 3047 439
rect 3049 435 3053 439
rect 3055 435 3059 439
rect 3061 435 3065 439
rect 3067 435 3071 439
rect 3073 435 3077 439
rect 3079 435 3083 439
rect 3043 429 3047 433
rect 3049 429 3053 433
rect 3055 429 3059 433
rect 3061 429 3065 433
rect 3067 429 3071 433
rect 3073 429 3077 433
rect 3079 429 3083 433
rect 3043 423 3047 427
rect 3049 423 3053 427
rect 3055 423 3059 427
rect 3061 423 3065 427
rect 3067 423 3071 427
rect 3073 423 3077 427
rect 3079 423 3083 427
rect 3043 412 3047 421
rect 3049 412 3053 421
rect 3055 412 3059 421
rect 3061 412 3065 421
rect 3067 412 3071 421
rect 3073 412 3077 421
rect 3079 412 3083 421
rect 2909 402 2913 406
rect 2915 402 2919 406
rect 2921 402 2925 406
rect 2927 402 2931 406
rect 2933 402 2937 406
rect 2939 402 2943 406
rect 2945 402 2949 406
rect 2909 390 2913 394
rect 2915 390 2919 394
rect 2921 390 2925 394
rect 2927 390 2931 394
rect 2933 390 2937 394
rect 2939 390 2943 394
rect 2945 390 2949 394
rect 2915 378 2919 382
rect 2921 378 2925 382
rect 2927 378 2931 382
rect 2933 378 2937 382
rect 2939 378 2943 382
rect 2945 378 2949 382
rect 2999 402 3003 406
rect 3005 402 3009 406
rect 3011 402 3015 406
rect 3017 402 3021 406
rect 3023 402 3027 406
rect 3029 402 3033 406
rect 3035 402 3039 406
rect 2999 390 3003 394
rect 3005 390 3009 394
rect 3011 390 3015 394
rect 3017 390 3021 394
rect 3023 390 3027 394
rect 3029 390 3033 394
rect 3035 390 3039 394
rect 2999 378 3003 382
rect 3005 378 3009 382
rect 3011 378 3015 382
rect 3017 378 3021 382
rect 3023 378 3027 382
rect 3029 378 3033 382
rect 3339 509 3343 513
rect 3345 509 3349 513
rect 3351 509 3355 513
rect 3357 509 3361 513
rect 3363 509 3367 513
rect 3369 509 3373 513
rect 3375 509 3379 513
rect 3339 441 3343 450
rect 3345 441 3349 450
rect 3351 441 3355 450
rect 3357 441 3361 450
rect 3363 441 3367 450
rect 3369 441 3373 450
rect 3375 441 3379 450
rect 3339 435 3343 439
rect 3345 435 3349 439
rect 3351 435 3355 439
rect 3357 435 3361 439
rect 3363 435 3367 439
rect 3369 435 3373 439
rect 3375 435 3379 439
rect 3339 429 3343 433
rect 3345 429 3349 433
rect 3351 429 3355 433
rect 3357 429 3361 433
rect 3363 429 3367 433
rect 3369 429 3373 433
rect 3375 429 3379 433
rect 3339 423 3343 427
rect 3345 423 3349 427
rect 3351 423 3355 427
rect 3357 423 3361 427
rect 3363 423 3367 427
rect 3369 423 3373 427
rect 3375 423 3379 427
rect 3339 412 3343 421
rect 3345 412 3349 421
rect 3351 412 3355 421
rect 3357 412 3361 421
rect 3363 412 3367 421
rect 3369 412 3373 421
rect 3375 412 3379 421
rect 3383 509 3387 513
rect 3389 509 3393 513
rect 3395 509 3399 513
rect 3401 509 3405 513
rect 3407 509 3411 513
rect 3413 509 3417 513
rect 3419 509 3423 513
rect 3389 495 3393 499
rect 3395 495 3399 499
rect 3401 495 3405 499
rect 3407 495 3411 499
rect 3413 495 3417 499
rect 3419 495 3423 499
rect 3383 483 3387 487
rect 3389 483 3393 487
rect 3395 483 3399 487
rect 3401 483 3405 487
rect 3407 483 3411 487
rect 3413 483 3417 487
rect 3419 483 3423 487
rect 3383 477 3387 481
rect 3389 477 3393 481
rect 3395 477 3399 481
rect 3401 477 3405 481
rect 3407 477 3411 481
rect 3413 477 3417 481
rect 3419 477 3423 481
rect 3383 465 3387 469
rect 3389 465 3393 469
rect 3395 465 3399 469
rect 3401 465 3405 469
rect 3407 465 3411 469
rect 3413 465 3417 469
rect 3419 465 3423 469
rect 3427 509 3436 513
rect 3422 456 3426 460
rect 3432 456 3436 460
rect 3460 509 3469 513
rect 3473 509 3477 513
rect 3479 509 3483 513
rect 3485 509 3489 513
rect 3491 509 3495 513
rect 3497 509 3501 513
rect 3503 509 3507 513
rect 3509 509 3513 513
rect 3473 495 3477 499
rect 3479 495 3483 499
rect 3485 495 3489 499
rect 3491 495 3495 499
rect 3497 495 3501 499
rect 3503 495 3507 499
rect 3473 483 3477 487
rect 3479 483 3483 487
rect 3485 483 3489 487
rect 3491 483 3495 487
rect 3497 483 3501 487
rect 3503 483 3507 487
rect 3509 483 3513 487
rect 3473 477 3477 481
rect 3479 477 3483 481
rect 3485 477 3489 481
rect 3491 477 3495 481
rect 3497 477 3501 481
rect 3503 477 3507 481
rect 3509 477 3513 481
rect 3473 465 3477 469
rect 3479 465 3483 469
rect 3485 465 3489 469
rect 3491 465 3495 469
rect 3497 465 3501 469
rect 3503 465 3507 469
rect 3509 465 3513 469
rect 3460 456 3464 460
rect 3470 456 3474 460
rect 3517 509 3521 513
rect 3523 509 3527 513
rect 3529 509 3533 513
rect 3535 509 3539 513
rect 3541 509 3545 513
rect 3547 509 3551 513
rect 3553 509 3557 513
rect 3517 441 3521 450
rect 3523 441 3527 450
rect 3529 441 3533 450
rect 3535 441 3539 450
rect 3541 441 3545 450
rect 3547 441 3551 450
rect 3553 441 3557 450
rect 3517 435 3521 439
rect 3523 435 3527 439
rect 3529 435 3533 439
rect 3535 435 3539 439
rect 3541 435 3545 439
rect 3547 435 3551 439
rect 3553 435 3557 439
rect 3517 429 3521 433
rect 3523 429 3527 433
rect 3529 429 3533 433
rect 3535 429 3539 433
rect 3541 429 3545 433
rect 3547 429 3551 433
rect 3553 429 3557 433
rect 3517 423 3521 427
rect 3523 423 3527 427
rect 3529 423 3533 427
rect 3535 423 3539 427
rect 3541 423 3545 427
rect 3547 423 3551 427
rect 3553 423 3557 427
rect 3517 412 3521 421
rect 3523 412 3527 421
rect 3529 412 3533 421
rect 3535 412 3539 421
rect 3541 412 3545 421
rect 3547 412 3551 421
rect 3553 412 3557 421
rect 3383 402 3387 406
rect 3389 402 3393 406
rect 3395 402 3399 406
rect 3401 402 3405 406
rect 3407 402 3411 406
rect 3413 402 3417 406
rect 3419 402 3423 406
rect 3383 390 3387 394
rect 3389 390 3393 394
rect 3395 390 3399 394
rect 3401 390 3405 394
rect 3407 390 3411 394
rect 3413 390 3417 394
rect 3419 390 3423 394
rect 3389 378 3393 382
rect 3395 378 3399 382
rect 3401 378 3405 382
rect 3407 378 3411 382
rect 3413 378 3417 382
rect 3419 378 3423 382
rect 3473 402 3477 406
rect 3479 402 3483 406
rect 3485 402 3489 406
rect 3491 402 3495 406
rect 3497 402 3501 406
rect 3503 402 3507 406
rect 3509 402 3513 406
rect 3473 390 3477 394
rect 3479 390 3483 394
rect 3485 390 3489 394
rect 3491 390 3495 394
rect 3497 390 3501 394
rect 3503 390 3507 394
rect 3509 390 3513 394
rect 3473 378 3477 382
rect 3479 378 3483 382
rect 3485 378 3489 382
rect 3491 378 3495 382
rect 3497 378 3501 382
rect 3503 378 3507 382
rect 3813 509 3817 513
rect 3819 509 3823 513
rect 3825 509 3829 513
rect 3831 509 3835 513
rect 3837 509 3841 513
rect 3843 509 3847 513
rect 3849 509 3853 513
rect 3813 441 3817 450
rect 3819 441 3823 450
rect 3825 441 3829 450
rect 3831 441 3835 450
rect 3837 441 3841 450
rect 3843 441 3847 450
rect 3849 441 3853 450
rect 3813 435 3817 439
rect 3819 435 3823 439
rect 3825 435 3829 439
rect 3831 435 3835 439
rect 3837 435 3841 439
rect 3843 435 3847 439
rect 3849 435 3853 439
rect 3813 429 3817 433
rect 3819 429 3823 433
rect 3825 429 3829 433
rect 3831 429 3835 433
rect 3837 429 3841 433
rect 3843 429 3847 433
rect 3849 429 3853 433
rect 3813 423 3817 427
rect 3819 423 3823 427
rect 3825 423 3829 427
rect 3831 423 3835 427
rect 3837 423 3841 427
rect 3843 423 3847 427
rect 3849 423 3853 427
rect 3813 412 3817 421
rect 3819 412 3823 421
rect 3825 412 3829 421
rect 3831 412 3835 421
rect 3837 412 3841 421
rect 3843 412 3847 421
rect 3849 412 3853 421
rect 3857 509 3861 513
rect 3863 509 3867 513
rect 3869 509 3873 513
rect 3875 509 3879 513
rect 3881 509 3885 513
rect 3887 509 3891 513
rect 3893 509 3897 513
rect 3863 495 3867 499
rect 3869 495 3873 499
rect 3875 495 3879 499
rect 3881 495 3885 499
rect 3887 495 3891 499
rect 3893 495 3897 499
rect 3857 483 3861 487
rect 3863 483 3867 487
rect 3869 483 3873 487
rect 3875 483 3879 487
rect 3881 483 3885 487
rect 3887 483 3891 487
rect 3893 483 3897 487
rect 3857 477 3861 481
rect 3863 477 3867 481
rect 3869 477 3873 481
rect 3875 477 3879 481
rect 3881 477 3885 481
rect 3887 477 3891 481
rect 3893 477 3897 481
rect 3857 465 3861 469
rect 3863 465 3867 469
rect 3869 465 3873 469
rect 3875 465 3879 469
rect 3881 465 3885 469
rect 3887 465 3891 469
rect 3893 465 3897 469
rect 3901 509 3910 513
rect 3896 456 3900 460
rect 3906 456 3910 460
rect 3934 509 3943 513
rect 3947 509 3951 513
rect 3953 509 3957 513
rect 3959 509 3963 513
rect 3965 509 3969 513
rect 3971 509 3975 513
rect 3977 509 3981 513
rect 3983 509 3987 513
rect 3947 495 3951 499
rect 3953 495 3957 499
rect 3959 495 3963 499
rect 3965 495 3969 499
rect 3971 495 3975 499
rect 3977 495 3981 499
rect 3947 483 3951 487
rect 3953 483 3957 487
rect 3959 483 3963 487
rect 3965 483 3969 487
rect 3971 483 3975 487
rect 3977 483 3981 487
rect 3983 483 3987 487
rect 3947 477 3951 481
rect 3953 477 3957 481
rect 3959 477 3963 481
rect 3965 477 3969 481
rect 3971 477 3975 481
rect 3977 477 3981 481
rect 3983 477 3987 481
rect 3947 465 3951 469
rect 3953 465 3957 469
rect 3959 465 3963 469
rect 3965 465 3969 469
rect 3971 465 3975 469
rect 3977 465 3981 469
rect 3983 465 3987 469
rect 3934 456 3938 460
rect 3944 456 3948 460
rect 3991 509 3995 513
rect 3997 509 4001 513
rect 4003 509 4007 513
rect 4009 509 4013 513
rect 4015 509 4019 513
rect 4021 509 4025 513
rect 4027 509 4031 513
rect 3991 441 3995 450
rect 3997 441 4001 450
rect 4003 441 4007 450
rect 4009 441 4013 450
rect 4015 441 4019 450
rect 4021 441 4025 450
rect 4027 441 4031 450
rect 3991 435 3995 439
rect 3997 435 4001 439
rect 4003 435 4007 439
rect 4009 435 4013 439
rect 4015 435 4019 439
rect 4021 435 4025 439
rect 4027 435 4031 439
rect 3991 429 3995 433
rect 3997 429 4001 433
rect 4003 429 4007 433
rect 4009 429 4013 433
rect 4015 429 4019 433
rect 4021 429 4025 433
rect 4027 429 4031 433
rect 3991 423 3995 427
rect 3997 423 4001 427
rect 4003 423 4007 427
rect 4009 423 4013 427
rect 4015 423 4019 427
rect 4021 423 4025 427
rect 4027 423 4031 427
rect 3991 412 3995 421
rect 3997 412 4001 421
rect 4003 412 4007 421
rect 4009 412 4013 421
rect 4015 412 4019 421
rect 4021 412 4025 421
rect 4027 412 4031 421
rect 3857 402 3861 406
rect 3863 402 3867 406
rect 3869 402 3873 406
rect 3875 402 3879 406
rect 3881 402 3885 406
rect 3887 402 3891 406
rect 3893 402 3897 406
rect 3857 390 3861 394
rect 3863 390 3867 394
rect 3869 390 3873 394
rect 3875 390 3879 394
rect 3881 390 3885 394
rect 3887 390 3891 394
rect 3893 390 3897 394
rect 3863 378 3867 382
rect 3869 378 3873 382
rect 3875 378 3879 382
rect 3881 378 3885 382
rect 3887 378 3891 382
rect 3893 378 3897 382
rect 3947 402 3951 406
rect 3953 402 3957 406
rect 3959 402 3963 406
rect 3965 402 3969 406
rect 3971 402 3975 406
rect 3977 402 3981 406
rect 3983 402 3987 406
rect 3947 390 3951 394
rect 3953 390 3957 394
rect 3959 390 3963 394
rect 3965 390 3969 394
rect 3971 390 3975 394
rect 3977 390 3981 394
rect 3983 390 3987 394
rect 3947 378 3951 382
rect 3953 378 3957 382
rect 3959 378 3963 382
rect 3965 378 3969 382
rect 3971 378 3975 382
rect 3977 378 3981 382
rect 4287 509 4291 513
rect 4293 509 4297 513
rect 4299 509 4303 513
rect 4305 509 4309 513
rect 4311 509 4315 513
rect 4317 509 4321 513
rect 4323 509 4327 513
rect 4287 441 4291 450
rect 4293 441 4297 450
rect 4299 441 4303 450
rect 4305 441 4309 450
rect 4311 441 4315 450
rect 4317 441 4321 450
rect 4323 441 4327 450
rect 4287 435 4291 439
rect 4293 435 4297 439
rect 4299 435 4303 439
rect 4305 435 4309 439
rect 4311 435 4315 439
rect 4317 435 4321 439
rect 4323 435 4327 439
rect 4287 429 4291 433
rect 4293 429 4297 433
rect 4299 429 4303 433
rect 4305 429 4309 433
rect 4311 429 4315 433
rect 4317 429 4321 433
rect 4323 429 4327 433
rect 4287 423 4291 427
rect 4293 423 4297 427
rect 4299 423 4303 427
rect 4305 423 4309 427
rect 4311 423 4315 427
rect 4317 423 4321 427
rect 4323 423 4327 427
rect 4287 412 4291 421
rect 4293 412 4297 421
rect 4299 412 4303 421
rect 4305 412 4309 421
rect 4311 412 4315 421
rect 4317 412 4321 421
rect 4323 412 4327 421
rect 4331 509 4335 513
rect 4337 509 4341 513
rect 4343 509 4347 513
rect 4349 509 4353 513
rect 4355 509 4359 513
rect 4361 509 4365 513
rect 4367 509 4371 513
rect 4337 495 4341 499
rect 4343 495 4347 499
rect 4349 495 4353 499
rect 4355 495 4359 499
rect 4361 495 4365 499
rect 4367 495 4371 499
rect 4331 483 4335 487
rect 4337 483 4341 487
rect 4343 483 4347 487
rect 4349 483 4353 487
rect 4355 483 4359 487
rect 4361 483 4365 487
rect 4367 483 4371 487
rect 4331 477 4335 481
rect 4337 477 4341 481
rect 4343 477 4347 481
rect 4349 477 4353 481
rect 4355 477 4359 481
rect 4361 477 4365 481
rect 4367 477 4371 481
rect 4331 465 4335 469
rect 4337 465 4341 469
rect 4343 465 4347 469
rect 4349 465 4353 469
rect 4355 465 4359 469
rect 4361 465 4365 469
rect 4367 465 4371 469
rect 4375 509 4384 513
rect 4370 456 4374 460
rect 4380 456 4384 460
rect 4408 509 4417 513
rect 4421 509 4425 513
rect 4427 509 4431 513
rect 4433 509 4437 513
rect 4439 509 4443 513
rect 4445 509 4449 513
rect 4451 509 4455 513
rect 4457 509 4461 513
rect 4421 495 4425 499
rect 4427 495 4431 499
rect 4433 495 4437 499
rect 4439 495 4443 499
rect 4445 495 4449 499
rect 4451 495 4455 499
rect 4457 495 4461 499
rect 4421 483 4425 487
rect 4427 483 4431 487
rect 4433 483 4437 487
rect 4439 483 4443 487
rect 4445 483 4449 487
rect 4451 483 4455 487
rect 4457 483 4461 487
rect 4421 477 4425 481
rect 4427 477 4431 481
rect 4433 477 4437 481
rect 4439 477 4443 481
rect 4445 477 4449 481
rect 4451 477 4455 481
rect 4457 477 4461 481
rect 4421 465 4425 469
rect 4427 465 4431 469
rect 4433 465 4437 469
rect 4439 465 4443 469
rect 4445 465 4449 469
rect 4451 465 4455 469
rect 4457 465 4461 469
rect 4408 456 4412 460
rect 4418 456 4422 460
rect 4465 441 4469 450
rect 4471 441 4475 450
rect 4477 441 4481 450
rect 4483 441 4487 450
rect 4489 441 4493 450
rect 4495 441 4499 450
rect 4501 441 4505 450
rect 4465 435 4469 439
rect 4471 435 4475 439
rect 4477 435 4481 439
rect 4483 435 4487 439
rect 4489 435 4493 439
rect 4495 435 4499 439
rect 4501 435 4505 439
rect 4465 429 4469 433
rect 4471 429 4475 433
rect 4477 429 4481 433
rect 4483 429 4487 433
rect 4489 429 4493 433
rect 4495 429 4499 433
rect 4501 429 4505 433
rect 4465 423 4469 427
rect 4471 423 4475 427
rect 4477 423 4481 427
rect 4483 423 4487 427
rect 4489 423 4493 427
rect 4495 423 4499 427
rect 4501 423 4505 427
rect 4465 412 4469 421
rect 4471 412 4475 421
rect 4477 412 4481 421
rect 4483 412 4487 421
rect 4489 412 4493 421
rect 4495 412 4499 421
rect 4501 412 4505 421
rect 4331 402 4335 406
rect 4337 402 4341 406
rect 4343 402 4347 406
rect 4349 402 4353 406
rect 4355 402 4359 406
rect 4361 402 4365 406
rect 4367 402 4371 406
rect 4331 390 4335 394
rect 4337 390 4341 394
rect 4343 390 4347 394
rect 4349 390 4353 394
rect 4355 390 4359 394
rect 4361 390 4365 394
rect 4367 390 4371 394
rect 4337 378 4341 382
rect 4343 378 4347 382
rect 4349 378 4353 382
rect 4355 378 4359 382
rect 4361 378 4365 382
rect 4367 378 4371 382
rect 4421 402 4425 406
rect 4427 402 4431 406
rect 4433 402 4437 406
rect 4439 402 4443 406
rect 4445 402 4449 406
rect 4451 402 4455 406
rect 4457 402 4461 406
rect 4421 390 4425 394
rect 4427 390 4431 394
rect 4433 390 4437 394
rect 4439 390 4443 394
rect 4445 390 4449 394
rect 4451 390 4455 394
rect 4457 390 4461 394
rect 4421 378 4425 382
rect 4427 378 4431 382
rect 4433 378 4437 382
rect 4439 378 4443 382
rect 4445 378 4449 382
rect 4451 378 4455 382
rect 327 255 331 259
rect 339 255 343 259
rect 351 255 355 259
rect 321 243 325 247
rect 333 243 337 247
rect 345 243 349 247
rect 327 231 331 235
rect 339 231 343 235
rect 351 231 355 235
rect 321 219 325 223
rect 333 219 337 223
rect 345 219 349 223
rect 4645 255 4649 259
rect 4657 255 4661 259
rect 4669 255 4673 259
rect 4651 243 4655 247
rect 4663 243 4667 247
rect 4675 243 4679 247
rect 4645 231 4649 235
rect 4657 231 4661 235
rect 4669 231 4673 235
rect 4651 219 4655 223
rect 4663 219 4667 223
rect 4675 219 4679 223
<< metal2 >>
rect 543 509 545 513
rect 549 509 551 513
rect 555 509 557 513
rect 561 509 563 513
rect 567 509 569 513
rect 573 509 575 513
rect 633 509 635 513
rect 639 509 641 513
rect 645 509 647 513
rect 651 509 653 513
rect 657 509 659 513
rect 663 509 665 513
rect 677 509 679 513
rect 683 509 685 513
rect 689 509 691 513
rect 695 509 697 513
rect 701 509 703 513
rect 707 509 709 513
rect 973 509 975 513
rect 979 509 981 513
rect 985 509 987 513
rect 991 509 993 513
rect 997 509 999 513
rect 1003 509 1005 513
rect 1017 509 1019 513
rect 1023 509 1025 513
rect 1029 509 1031 513
rect 1035 509 1037 513
rect 1041 509 1043 513
rect 1047 509 1049 513
rect 1107 509 1109 513
rect 1113 509 1115 513
rect 1119 509 1121 513
rect 1125 509 1127 513
rect 1131 509 1133 513
rect 1137 509 1139 513
rect 1151 509 1153 513
rect 1157 509 1159 513
rect 1163 509 1165 513
rect 1169 509 1171 513
rect 1175 509 1177 513
rect 1181 509 1183 513
rect 1447 509 1449 513
rect 1453 509 1455 513
rect 1459 509 1461 513
rect 1465 509 1467 513
rect 1471 509 1473 513
rect 1477 509 1479 513
rect 1491 509 1493 513
rect 1497 509 1499 513
rect 1503 509 1505 513
rect 1509 509 1511 513
rect 1515 509 1517 513
rect 1521 509 1523 513
rect 1581 509 1583 513
rect 1587 509 1589 513
rect 1593 509 1595 513
rect 1599 509 1601 513
rect 1605 509 1607 513
rect 1611 509 1613 513
rect 1625 509 1627 513
rect 1631 509 1633 513
rect 1637 509 1639 513
rect 1643 509 1645 513
rect 1649 509 1651 513
rect 1655 509 1657 513
rect 1921 509 1923 513
rect 1927 509 1929 513
rect 1933 509 1935 513
rect 1939 509 1941 513
rect 1945 509 1947 513
rect 1951 509 1953 513
rect 1965 509 1967 513
rect 1971 509 1973 513
rect 1977 509 1979 513
rect 1983 509 1985 513
rect 1989 509 1991 513
rect 1995 509 1997 513
rect 2055 509 2057 513
rect 2061 509 2063 513
rect 2067 509 2069 513
rect 2073 509 2075 513
rect 2079 509 2081 513
rect 2085 509 2087 513
rect 2099 509 2101 513
rect 2105 509 2107 513
rect 2111 509 2113 513
rect 2117 509 2119 513
rect 2123 509 2125 513
rect 2129 509 2131 513
rect 2395 509 2397 513
rect 2401 509 2403 513
rect 2407 509 2409 513
rect 2413 509 2415 513
rect 2419 509 2421 513
rect 2425 509 2427 513
rect 2439 509 2441 513
rect 2445 509 2447 513
rect 2451 509 2453 513
rect 2457 509 2459 513
rect 2463 509 2465 513
rect 2469 509 2471 513
rect 2529 509 2531 513
rect 2535 509 2537 513
rect 2541 509 2543 513
rect 2547 509 2549 513
rect 2553 509 2555 513
rect 2559 509 2561 513
rect 2573 509 2575 513
rect 2579 509 2581 513
rect 2585 509 2587 513
rect 2591 509 2593 513
rect 2597 509 2599 513
rect 2603 509 2605 513
rect 2869 509 2871 513
rect 2875 509 2877 513
rect 2881 509 2883 513
rect 2887 509 2889 513
rect 2893 509 2895 513
rect 2899 509 2901 513
rect 2913 509 2915 513
rect 2919 509 2921 513
rect 2925 509 2927 513
rect 2931 509 2933 513
rect 2937 509 2939 513
rect 2943 509 2945 513
rect 3003 509 3005 513
rect 3009 509 3011 513
rect 3015 509 3017 513
rect 3021 509 3023 513
rect 3027 509 3029 513
rect 3033 509 3035 513
rect 3047 509 3049 513
rect 3053 509 3055 513
rect 3059 509 3061 513
rect 3065 509 3067 513
rect 3071 509 3073 513
rect 3077 509 3079 513
rect 3343 509 3345 513
rect 3349 509 3351 513
rect 3355 509 3357 513
rect 3361 509 3363 513
rect 3367 509 3369 513
rect 3373 509 3375 513
rect 3387 509 3389 513
rect 3393 509 3395 513
rect 3399 509 3401 513
rect 3405 509 3407 513
rect 3411 509 3413 513
rect 3417 509 3419 513
rect 3477 509 3479 513
rect 3483 509 3485 513
rect 3489 509 3491 513
rect 3495 509 3497 513
rect 3501 509 3503 513
rect 3507 509 3509 513
rect 3521 509 3523 513
rect 3527 509 3529 513
rect 3533 509 3535 513
rect 3539 509 3541 513
rect 3545 509 3547 513
rect 3551 509 3553 513
rect 3817 509 3819 513
rect 3823 509 3825 513
rect 3829 509 3831 513
rect 3835 509 3837 513
rect 3841 509 3843 513
rect 3847 509 3849 513
rect 3861 509 3863 513
rect 3867 509 3869 513
rect 3873 509 3875 513
rect 3879 509 3881 513
rect 3885 509 3887 513
rect 3891 509 3893 513
rect 3951 509 3953 513
rect 3957 509 3959 513
rect 3963 509 3965 513
rect 3969 509 3971 513
rect 3975 509 3977 513
rect 3981 509 3983 513
rect 3995 509 3997 513
rect 4001 509 4003 513
rect 4007 509 4009 513
rect 4013 509 4015 513
rect 4019 509 4021 513
rect 4025 509 4027 513
rect 4291 509 4293 513
rect 4297 509 4299 513
rect 4303 509 4305 513
rect 4309 509 4311 513
rect 4315 509 4317 513
rect 4321 509 4323 513
rect 4335 509 4337 513
rect 4341 509 4343 513
rect 4347 509 4349 513
rect 4353 509 4355 513
rect 4359 509 4361 513
rect 4365 509 4367 513
rect 4425 509 4427 513
rect 4431 509 4433 513
rect 4437 509 4439 513
rect 4443 509 4445 513
rect 4449 509 4451 513
rect 4455 509 4457 513
rect 539 505 579 509
rect 629 505 669 509
rect 1013 505 1053 509
rect 1103 505 1143 509
rect 1487 505 1527 509
rect 1577 505 1617 509
rect 1961 505 2001 509
rect 2051 505 2091 509
rect 2435 505 2475 509
rect 2525 505 2565 509
rect 2909 505 2949 509
rect 2999 505 3039 509
rect 3383 505 3423 509
rect 3473 505 3513 509
rect 3857 505 3897 509
rect 3947 505 3987 509
rect 4331 505 4371 509
rect 4421 505 4461 509
rect 465 499 4535 505
rect 465 496 539 499
rect 465 467 467 496
rect 531 495 539 496
rect 543 495 545 499
rect 549 495 551 499
rect 555 495 557 499
rect 561 495 563 499
rect 567 495 569 499
rect 573 495 575 499
rect 579 495 629 499
rect 633 495 635 499
rect 639 495 641 499
rect 645 495 647 499
rect 651 495 653 499
rect 657 495 659 499
rect 663 495 1019 499
rect 1023 495 1025 499
rect 1029 495 1031 499
rect 1035 495 1037 499
rect 1041 495 1043 499
rect 1047 495 1049 499
rect 1053 495 1103 499
rect 1107 495 1109 499
rect 1113 495 1115 499
rect 1119 495 1121 499
rect 1125 495 1127 499
rect 1131 495 1133 499
rect 1137 495 1493 499
rect 1497 495 1499 499
rect 1503 495 1505 499
rect 1509 495 1511 499
rect 1515 495 1517 499
rect 1521 495 1523 499
rect 1527 495 1577 499
rect 1581 495 1583 499
rect 1587 495 1589 499
rect 1593 495 1595 499
rect 1599 495 1601 499
rect 1605 495 1607 499
rect 1611 495 1967 499
rect 1971 495 1973 499
rect 1977 495 1979 499
rect 1983 495 1985 499
rect 1989 495 1991 499
rect 1995 495 1997 499
rect 2001 495 2051 499
rect 2055 495 2057 499
rect 2061 495 2063 499
rect 2067 495 2069 499
rect 2073 495 2075 499
rect 2079 495 2081 499
rect 2085 495 2441 499
rect 2445 495 2447 499
rect 2451 495 2453 499
rect 2457 495 2459 499
rect 2463 495 2465 499
rect 2469 495 2471 499
rect 2475 495 2525 499
rect 2529 495 2531 499
rect 2535 495 2537 499
rect 2541 495 2543 499
rect 2547 495 2549 499
rect 2553 495 2555 499
rect 2559 495 2915 499
rect 2919 495 2921 499
rect 2925 495 2927 499
rect 2931 495 2933 499
rect 2937 495 2939 499
rect 2943 495 2945 499
rect 2949 495 2999 499
rect 3003 495 3005 499
rect 3009 495 3011 499
rect 3015 495 3017 499
rect 3021 495 3023 499
rect 3027 495 3029 499
rect 3033 495 3389 499
rect 3393 495 3395 499
rect 3399 495 3401 499
rect 3405 495 3407 499
rect 3411 495 3413 499
rect 3417 495 3419 499
rect 3423 495 3473 499
rect 3477 495 3479 499
rect 3483 495 3485 499
rect 3489 495 3491 499
rect 3495 495 3497 499
rect 3501 495 3503 499
rect 3507 495 3863 499
rect 3867 495 3869 499
rect 3873 495 3875 499
rect 3879 495 3881 499
rect 3885 495 3887 499
rect 3891 495 3893 499
rect 3897 495 3947 499
rect 3951 495 3953 499
rect 3957 495 3959 499
rect 3963 495 3965 499
rect 3969 495 3971 499
rect 3975 495 3977 499
rect 3981 495 4337 499
rect 4341 495 4343 499
rect 4347 495 4349 499
rect 4353 495 4355 499
rect 4359 495 4361 499
rect 4365 495 4367 499
rect 4371 495 4421 499
rect 4425 495 4427 499
rect 4431 495 4433 499
rect 4437 495 4439 499
rect 4443 495 4445 499
rect 4449 495 4451 499
rect 4455 495 4457 499
rect 4461 495 4535 499
rect 531 487 4535 495
rect 531 483 539 487
rect 543 483 545 487
rect 549 483 551 487
rect 555 483 557 487
rect 561 483 563 487
rect 567 483 569 487
rect 573 483 575 487
rect 579 483 629 487
rect 633 483 635 487
rect 639 483 641 487
rect 645 483 647 487
rect 651 483 653 487
rect 657 483 659 487
rect 663 483 665 487
rect 669 483 1013 487
rect 1017 483 1019 487
rect 1023 483 1025 487
rect 1029 483 1031 487
rect 1035 483 1037 487
rect 1041 483 1043 487
rect 1047 483 1049 487
rect 1053 483 1103 487
rect 1107 483 1109 487
rect 1113 483 1115 487
rect 1119 483 1121 487
rect 1125 483 1127 487
rect 1131 483 1133 487
rect 1137 483 1139 487
rect 1143 483 1487 487
rect 1491 483 1493 487
rect 1497 483 1499 487
rect 1503 483 1505 487
rect 1509 483 1511 487
rect 1515 483 1517 487
rect 1521 483 1523 487
rect 1527 483 1577 487
rect 1581 483 1583 487
rect 1587 483 1589 487
rect 1593 483 1595 487
rect 1599 483 1601 487
rect 1605 483 1607 487
rect 1611 483 1613 487
rect 1617 483 1961 487
rect 1965 483 1967 487
rect 1971 483 1973 487
rect 1977 483 1979 487
rect 1983 483 1985 487
rect 1989 483 1991 487
rect 1995 483 1997 487
rect 2001 483 2051 487
rect 2055 483 2057 487
rect 2061 483 2063 487
rect 2067 483 2069 487
rect 2073 483 2075 487
rect 2079 483 2081 487
rect 2085 483 2087 487
rect 2091 483 2435 487
rect 2439 483 2441 487
rect 2445 483 2447 487
rect 2451 483 2453 487
rect 2457 483 2459 487
rect 2463 483 2465 487
rect 2469 483 2471 487
rect 2475 483 2525 487
rect 2529 483 2531 487
rect 2535 483 2537 487
rect 2541 483 2543 487
rect 2547 483 2549 487
rect 2553 483 2555 487
rect 2559 483 2561 487
rect 2565 483 2909 487
rect 2913 483 2915 487
rect 2919 483 2921 487
rect 2925 483 2927 487
rect 2931 483 2933 487
rect 2937 483 2939 487
rect 2943 483 2945 487
rect 2949 483 2999 487
rect 3003 483 3005 487
rect 3009 483 3011 487
rect 3015 483 3017 487
rect 3021 483 3023 487
rect 3027 483 3029 487
rect 3033 483 3035 487
rect 3039 483 3383 487
rect 3387 483 3389 487
rect 3393 483 3395 487
rect 3399 483 3401 487
rect 3405 483 3407 487
rect 3411 483 3413 487
rect 3417 483 3419 487
rect 3423 483 3473 487
rect 3477 483 3479 487
rect 3483 483 3485 487
rect 3489 483 3491 487
rect 3495 483 3497 487
rect 3501 483 3503 487
rect 3507 483 3509 487
rect 3513 483 3857 487
rect 3861 483 3863 487
rect 3867 483 3869 487
rect 3873 483 3875 487
rect 3879 483 3881 487
rect 3885 483 3887 487
rect 3891 483 3893 487
rect 3897 483 3947 487
rect 3951 483 3953 487
rect 3957 483 3959 487
rect 3963 483 3965 487
rect 3969 483 3971 487
rect 3975 483 3977 487
rect 3981 483 3983 487
rect 3987 483 4331 487
rect 4335 483 4337 487
rect 4341 483 4343 487
rect 4347 483 4349 487
rect 4353 483 4355 487
rect 4359 483 4361 487
rect 4365 483 4367 487
rect 4371 483 4421 487
rect 4425 483 4427 487
rect 4431 483 4433 487
rect 4437 483 4439 487
rect 4443 483 4445 487
rect 4449 483 4451 487
rect 4455 483 4457 487
rect 4461 483 4535 487
rect 531 481 4535 483
rect 531 477 539 481
rect 543 477 545 481
rect 549 477 551 481
rect 555 477 557 481
rect 561 477 563 481
rect 567 477 569 481
rect 573 477 575 481
rect 579 477 629 481
rect 633 477 635 481
rect 639 477 641 481
rect 645 477 647 481
rect 651 477 653 481
rect 657 477 659 481
rect 663 477 665 481
rect 669 477 1013 481
rect 1017 477 1019 481
rect 1023 477 1025 481
rect 1029 477 1031 481
rect 1035 477 1037 481
rect 1041 477 1043 481
rect 1047 477 1049 481
rect 1053 477 1103 481
rect 1107 477 1109 481
rect 1113 477 1115 481
rect 1119 477 1121 481
rect 1125 477 1127 481
rect 1131 477 1133 481
rect 1137 477 1139 481
rect 1143 477 1487 481
rect 1491 477 1493 481
rect 1497 477 1499 481
rect 1503 477 1505 481
rect 1509 477 1511 481
rect 1515 477 1517 481
rect 1521 477 1523 481
rect 1527 477 1577 481
rect 1581 477 1583 481
rect 1587 477 1589 481
rect 1593 477 1595 481
rect 1599 477 1601 481
rect 1605 477 1607 481
rect 1611 477 1613 481
rect 1617 477 1961 481
rect 1965 477 1967 481
rect 1971 477 1973 481
rect 1977 477 1979 481
rect 1983 477 1985 481
rect 1989 477 1991 481
rect 1995 477 1997 481
rect 2001 477 2051 481
rect 2055 477 2057 481
rect 2061 477 2063 481
rect 2067 477 2069 481
rect 2073 477 2075 481
rect 2079 477 2081 481
rect 2085 477 2087 481
rect 2091 477 2435 481
rect 2439 477 2441 481
rect 2445 477 2447 481
rect 2451 477 2453 481
rect 2457 477 2459 481
rect 2463 477 2465 481
rect 2469 477 2471 481
rect 2475 477 2525 481
rect 2529 477 2531 481
rect 2535 477 2537 481
rect 2541 477 2543 481
rect 2547 477 2549 481
rect 2553 477 2555 481
rect 2559 477 2561 481
rect 2565 477 2909 481
rect 2913 477 2915 481
rect 2919 477 2921 481
rect 2925 477 2927 481
rect 2931 477 2933 481
rect 2937 477 2939 481
rect 2943 477 2945 481
rect 2949 477 2999 481
rect 3003 477 3005 481
rect 3009 477 3011 481
rect 3015 477 3017 481
rect 3021 477 3023 481
rect 3027 477 3029 481
rect 3033 477 3035 481
rect 3039 477 3383 481
rect 3387 477 3389 481
rect 3393 477 3395 481
rect 3399 477 3401 481
rect 3405 477 3407 481
rect 3411 477 3413 481
rect 3417 477 3419 481
rect 3423 477 3473 481
rect 3477 477 3479 481
rect 3483 477 3485 481
rect 3489 477 3491 481
rect 3495 477 3497 481
rect 3501 477 3503 481
rect 3507 477 3509 481
rect 3513 477 3857 481
rect 3861 477 3863 481
rect 3867 477 3869 481
rect 3873 477 3875 481
rect 3879 477 3881 481
rect 3885 477 3887 481
rect 3891 477 3893 481
rect 3897 477 3947 481
rect 3951 477 3953 481
rect 3957 477 3959 481
rect 3963 477 3965 481
rect 3969 477 3971 481
rect 3975 477 3977 481
rect 3981 477 3983 481
rect 3987 477 4331 481
rect 4335 477 4337 481
rect 4341 477 4343 481
rect 4347 477 4349 481
rect 4353 477 4355 481
rect 4359 477 4361 481
rect 4365 477 4367 481
rect 4371 477 4421 481
rect 4425 477 4427 481
rect 4431 477 4433 481
rect 4437 477 4439 481
rect 4443 477 4445 481
rect 4449 477 4451 481
rect 4455 477 4457 481
rect 4461 477 4535 481
rect 531 470 4535 477
rect 531 467 539 470
rect 465 466 539 467
rect 543 466 545 470
rect 549 466 551 470
rect 555 466 557 470
rect 561 466 563 470
rect 567 466 569 470
rect 573 466 575 470
rect 579 466 629 470
rect 633 466 635 470
rect 639 466 641 470
rect 645 466 647 470
rect 651 466 653 470
rect 657 466 659 470
rect 663 466 665 470
rect 669 469 4535 470
rect 669 466 1013 469
rect 465 465 1013 466
rect 1017 465 1019 469
rect 1023 465 1025 469
rect 1029 465 1031 469
rect 1035 465 1037 469
rect 1041 465 1043 469
rect 1047 465 1049 469
rect 1053 465 1103 469
rect 1107 465 1109 469
rect 1113 465 1115 469
rect 1119 465 1121 469
rect 1125 465 1127 469
rect 1131 465 1133 469
rect 1137 465 1139 469
rect 1143 465 1487 469
rect 1491 465 1493 469
rect 1497 465 1499 469
rect 1503 465 1505 469
rect 1509 465 1511 469
rect 1515 465 1517 469
rect 1521 465 1523 469
rect 1527 465 1577 469
rect 1581 465 1583 469
rect 1587 465 1589 469
rect 1593 465 1595 469
rect 1599 465 1601 469
rect 1605 465 1607 469
rect 1611 465 1613 469
rect 1617 465 1961 469
rect 1965 465 1967 469
rect 1971 465 1973 469
rect 1977 465 1979 469
rect 1983 465 1985 469
rect 1989 465 1991 469
rect 1995 465 1997 469
rect 2001 465 2051 469
rect 2055 465 2057 469
rect 2061 465 2063 469
rect 2067 465 2069 469
rect 2073 465 2075 469
rect 2079 465 2081 469
rect 2085 465 2087 469
rect 2091 465 2435 469
rect 2439 465 2441 469
rect 2445 465 2447 469
rect 2451 465 2453 469
rect 2457 465 2459 469
rect 2463 465 2465 469
rect 2469 465 2471 469
rect 2475 465 2525 469
rect 2529 465 2531 469
rect 2535 465 2537 469
rect 2541 465 2543 469
rect 2547 465 2549 469
rect 2553 465 2555 469
rect 2559 465 2561 469
rect 2565 465 2909 469
rect 2913 465 2915 469
rect 2919 465 2921 469
rect 2925 465 2927 469
rect 2931 465 2933 469
rect 2937 465 2939 469
rect 2943 465 2945 469
rect 2949 465 2999 469
rect 3003 465 3005 469
rect 3009 465 3011 469
rect 3015 465 3017 469
rect 3021 465 3023 469
rect 3027 465 3029 469
rect 3033 465 3035 469
rect 3039 465 3383 469
rect 3387 465 3389 469
rect 3393 465 3395 469
rect 3399 465 3401 469
rect 3405 465 3407 469
rect 3411 465 3413 469
rect 3417 465 3419 469
rect 3423 465 3473 469
rect 3477 465 3479 469
rect 3483 465 3485 469
rect 3489 465 3491 469
rect 3495 465 3497 469
rect 3501 465 3503 469
rect 3507 465 3509 469
rect 3513 465 3857 469
rect 3861 465 3863 469
rect 3867 465 3869 469
rect 3873 465 3875 469
rect 3879 465 3881 469
rect 3885 465 3887 469
rect 3891 465 3893 469
rect 3897 465 3947 469
rect 3951 465 3953 469
rect 3957 465 3959 469
rect 3963 465 3965 469
rect 3969 465 3971 469
rect 3975 465 3977 469
rect 3981 465 3983 469
rect 3987 465 4331 469
rect 4335 465 4337 469
rect 4341 465 4343 469
rect 4347 465 4349 469
rect 4353 465 4355 469
rect 4359 465 4361 469
rect 4365 465 4367 469
rect 4371 465 4421 469
rect 4425 465 4427 469
rect 4431 465 4433 469
rect 4437 465 4439 469
rect 4443 465 4445 469
rect 4449 465 4451 469
rect 4455 465 4457 469
rect 4461 465 4535 469
rect 455 460 4545 461
rect 455 456 578 460
rect 582 456 588 460
rect 592 456 616 460
rect 620 456 626 460
rect 630 456 1052 460
rect 1056 456 1062 460
rect 1066 456 1090 460
rect 1094 456 1100 460
rect 1104 456 1526 460
rect 1530 456 1536 460
rect 1540 456 1564 460
rect 1568 456 1574 460
rect 1578 456 2000 460
rect 2004 456 2010 460
rect 2014 456 2038 460
rect 2042 456 2048 460
rect 2052 456 2474 460
rect 2478 456 2484 460
rect 2488 456 2512 460
rect 2516 456 2522 460
rect 2526 456 2948 460
rect 2952 456 2958 460
rect 2962 456 2986 460
rect 2990 456 2996 460
rect 3000 456 3422 460
rect 3426 456 3432 460
rect 3436 456 3460 460
rect 3464 456 3470 460
rect 3474 456 3896 460
rect 3900 456 3906 460
rect 3910 456 3934 460
rect 3938 456 3944 460
rect 3948 456 4370 460
rect 4374 456 4380 460
rect 4384 456 4408 460
rect 4412 456 4418 460
rect 4422 456 4545 460
rect 455 455 4545 456
rect 411 450 4589 451
rect 411 441 495 450
rect 499 441 501 450
rect 505 441 507 450
rect 511 441 513 450
rect 517 441 519 450
rect 523 441 525 450
rect 529 441 531 450
rect 535 441 673 450
rect 677 441 679 450
rect 683 441 685 450
rect 689 441 691 450
rect 695 441 697 450
rect 701 441 703 450
rect 707 441 709 450
rect 713 441 969 450
rect 973 441 975 450
rect 979 441 981 450
rect 985 441 987 450
rect 991 441 993 450
rect 997 441 999 450
rect 1003 441 1005 450
rect 1009 441 1147 450
rect 1151 441 1153 450
rect 1157 441 1159 450
rect 1163 441 1165 450
rect 1169 441 1171 450
rect 1175 441 1177 450
rect 1181 441 1183 450
rect 1187 441 1443 450
rect 1447 441 1449 450
rect 1453 441 1455 450
rect 1459 441 1461 450
rect 1465 441 1467 450
rect 1471 441 1473 450
rect 1477 441 1479 450
rect 1483 441 1621 450
rect 1625 441 1627 450
rect 1631 441 1633 450
rect 1637 441 1639 450
rect 1643 441 1645 450
rect 1649 441 1651 450
rect 1655 441 1657 450
rect 1661 441 1917 450
rect 1921 441 1923 450
rect 1927 441 1929 450
rect 1933 441 1935 450
rect 1939 441 1941 450
rect 1945 441 1947 450
rect 1951 441 1953 450
rect 1957 441 2095 450
rect 2099 441 2101 450
rect 2105 441 2107 450
rect 2111 441 2113 450
rect 2117 441 2119 450
rect 2123 441 2125 450
rect 2129 441 2131 450
rect 2135 441 2391 450
rect 2395 441 2397 450
rect 2401 441 2403 450
rect 2407 441 2409 450
rect 2413 441 2415 450
rect 2419 441 2421 450
rect 2425 441 2427 450
rect 2431 441 2569 450
rect 2573 441 2575 450
rect 2579 441 2581 450
rect 2585 441 2587 450
rect 2591 441 2593 450
rect 2597 441 2599 450
rect 2603 441 2605 450
rect 2609 441 2865 450
rect 2869 441 2871 450
rect 2875 441 2877 450
rect 2881 441 2883 450
rect 2887 441 2889 450
rect 2893 441 2895 450
rect 2899 441 2901 450
rect 2905 441 3043 450
rect 3047 441 3049 450
rect 3053 441 3055 450
rect 3059 441 3061 450
rect 3065 441 3067 450
rect 3071 441 3073 450
rect 3077 441 3079 450
rect 3083 441 3339 450
rect 3343 441 3345 450
rect 3349 441 3351 450
rect 3355 441 3357 450
rect 3361 441 3363 450
rect 3367 441 3369 450
rect 3373 441 3375 450
rect 3379 441 3517 450
rect 3521 441 3523 450
rect 3527 441 3529 450
rect 3533 441 3535 450
rect 3539 441 3541 450
rect 3545 441 3547 450
rect 3551 441 3553 450
rect 3557 441 3813 450
rect 3817 441 3819 450
rect 3823 441 3825 450
rect 3829 441 3831 450
rect 3835 441 3837 450
rect 3841 441 3843 450
rect 3847 441 3849 450
rect 3853 441 3991 450
rect 3995 441 3997 450
rect 4001 441 4003 450
rect 4007 441 4009 450
rect 4013 441 4015 450
rect 4019 441 4021 450
rect 4025 441 4027 450
rect 4031 441 4287 450
rect 4291 441 4293 450
rect 4297 441 4299 450
rect 4303 441 4305 450
rect 4309 441 4311 450
rect 4315 441 4317 450
rect 4321 441 4323 450
rect 4327 441 4465 450
rect 4469 441 4471 450
rect 4475 441 4477 450
rect 4481 441 4483 450
rect 4487 441 4489 450
rect 4493 441 4495 450
rect 4499 441 4501 450
rect 4505 441 4589 450
rect 411 439 4589 441
rect 411 435 495 439
rect 499 435 501 439
rect 505 435 507 439
rect 511 435 513 439
rect 517 435 519 439
rect 523 435 525 439
rect 529 435 531 439
rect 535 435 673 439
rect 677 435 679 439
rect 683 435 685 439
rect 689 435 691 439
rect 695 435 697 439
rect 701 435 703 439
rect 707 435 709 439
rect 713 435 969 439
rect 973 435 975 439
rect 979 435 981 439
rect 985 435 987 439
rect 991 435 993 439
rect 997 435 999 439
rect 1003 435 1005 439
rect 1009 435 1147 439
rect 1151 435 1153 439
rect 1157 435 1159 439
rect 1163 435 1165 439
rect 1169 435 1171 439
rect 1175 435 1177 439
rect 1181 435 1183 439
rect 1187 435 1443 439
rect 1447 435 1449 439
rect 1453 435 1455 439
rect 1459 435 1461 439
rect 1465 435 1467 439
rect 1471 435 1473 439
rect 1477 435 1479 439
rect 1483 435 1621 439
rect 1625 435 1627 439
rect 1631 435 1633 439
rect 1637 435 1639 439
rect 1643 435 1645 439
rect 1649 435 1651 439
rect 1655 435 1657 439
rect 1661 435 1917 439
rect 1921 435 1923 439
rect 1927 435 1929 439
rect 1933 435 1935 439
rect 1939 435 1941 439
rect 1945 435 1947 439
rect 1951 435 1953 439
rect 1957 435 2095 439
rect 2099 435 2101 439
rect 2105 435 2107 439
rect 2111 435 2113 439
rect 2117 435 2119 439
rect 2123 435 2125 439
rect 2129 435 2131 439
rect 2135 435 2391 439
rect 2395 435 2397 439
rect 2401 435 2403 439
rect 2407 435 2409 439
rect 2413 435 2415 439
rect 2419 435 2421 439
rect 2425 435 2427 439
rect 2431 435 2569 439
rect 2573 435 2575 439
rect 2579 435 2581 439
rect 2585 435 2587 439
rect 2591 435 2593 439
rect 2597 435 2599 439
rect 2603 435 2605 439
rect 2609 435 2865 439
rect 2869 435 2871 439
rect 2875 435 2877 439
rect 2881 435 2883 439
rect 2887 435 2889 439
rect 2893 435 2895 439
rect 2899 435 2901 439
rect 2905 435 3043 439
rect 3047 435 3049 439
rect 3053 435 3055 439
rect 3059 435 3061 439
rect 3065 435 3067 439
rect 3071 435 3073 439
rect 3077 435 3079 439
rect 3083 435 3339 439
rect 3343 435 3345 439
rect 3349 435 3351 439
rect 3355 435 3357 439
rect 3361 435 3363 439
rect 3367 435 3369 439
rect 3373 435 3375 439
rect 3379 435 3517 439
rect 3521 435 3523 439
rect 3527 435 3529 439
rect 3533 435 3535 439
rect 3539 435 3541 439
rect 3545 435 3547 439
rect 3551 435 3553 439
rect 3557 435 3813 439
rect 3817 435 3819 439
rect 3823 435 3825 439
rect 3829 435 3831 439
rect 3835 435 3837 439
rect 3841 435 3843 439
rect 3847 435 3849 439
rect 3853 435 3991 439
rect 3995 435 3997 439
rect 4001 435 4003 439
rect 4007 435 4009 439
rect 4013 435 4015 439
rect 4019 435 4021 439
rect 4025 435 4027 439
rect 4031 435 4287 439
rect 4291 435 4293 439
rect 4297 435 4299 439
rect 4303 435 4305 439
rect 4309 435 4311 439
rect 4315 435 4317 439
rect 4321 435 4323 439
rect 4327 435 4465 439
rect 4469 435 4471 439
rect 4475 435 4477 439
rect 4481 435 4483 439
rect 4487 435 4489 439
rect 4493 435 4495 439
rect 4499 435 4501 439
rect 4505 435 4589 439
rect 411 433 4589 435
rect 411 429 495 433
rect 499 429 501 433
rect 505 429 507 433
rect 511 429 513 433
rect 517 429 519 433
rect 523 429 525 433
rect 529 429 531 433
rect 535 429 673 433
rect 677 429 679 433
rect 683 429 685 433
rect 689 429 691 433
rect 695 429 697 433
rect 701 429 703 433
rect 707 429 709 433
rect 713 429 969 433
rect 973 429 975 433
rect 979 429 981 433
rect 985 429 987 433
rect 991 429 993 433
rect 997 429 999 433
rect 1003 429 1005 433
rect 1009 429 1147 433
rect 1151 429 1153 433
rect 1157 429 1159 433
rect 1163 429 1165 433
rect 1169 429 1171 433
rect 1175 429 1177 433
rect 1181 429 1183 433
rect 1187 429 1443 433
rect 1447 429 1449 433
rect 1453 429 1455 433
rect 1459 429 1461 433
rect 1465 429 1467 433
rect 1471 429 1473 433
rect 1477 429 1479 433
rect 1483 429 1621 433
rect 1625 429 1627 433
rect 1631 429 1633 433
rect 1637 429 1639 433
rect 1643 429 1645 433
rect 1649 429 1651 433
rect 1655 429 1657 433
rect 1661 429 1917 433
rect 1921 429 1923 433
rect 1927 429 1929 433
rect 1933 429 1935 433
rect 1939 429 1941 433
rect 1945 429 1947 433
rect 1951 429 1953 433
rect 1957 429 2095 433
rect 2099 429 2101 433
rect 2105 429 2107 433
rect 2111 429 2113 433
rect 2117 429 2119 433
rect 2123 429 2125 433
rect 2129 429 2131 433
rect 2135 429 2391 433
rect 2395 429 2397 433
rect 2401 429 2403 433
rect 2407 429 2409 433
rect 2413 429 2415 433
rect 2419 429 2421 433
rect 2425 429 2427 433
rect 2431 429 2569 433
rect 2573 429 2575 433
rect 2579 429 2581 433
rect 2585 429 2587 433
rect 2591 429 2593 433
rect 2597 429 2599 433
rect 2603 429 2605 433
rect 2609 429 2865 433
rect 2869 429 2871 433
rect 2875 429 2877 433
rect 2881 429 2883 433
rect 2887 429 2889 433
rect 2893 429 2895 433
rect 2899 429 2901 433
rect 2905 429 3043 433
rect 3047 429 3049 433
rect 3053 429 3055 433
rect 3059 429 3061 433
rect 3065 429 3067 433
rect 3071 429 3073 433
rect 3077 429 3079 433
rect 3083 429 3339 433
rect 3343 429 3345 433
rect 3349 429 3351 433
rect 3355 429 3357 433
rect 3361 429 3363 433
rect 3367 429 3369 433
rect 3373 429 3375 433
rect 3379 429 3517 433
rect 3521 429 3523 433
rect 3527 429 3529 433
rect 3533 429 3535 433
rect 3539 429 3541 433
rect 3545 429 3547 433
rect 3551 429 3553 433
rect 3557 429 3813 433
rect 3817 429 3819 433
rect 3823 429 3825 433
rect 3829 429 3831 433
rect 3835 429 3837 433
rect 3841 429 3843 433
rect 3847 429 3849 433
rect 3853 429 3991 433
rect 3995 429 3997 433
rect 4001 429 4003 433
rect 4007 429 4009 433
rect 4013 429 4015 433
rect 4019 429 4021 433
rect 4025 429 4027 433
rect 4031 429 4287 433
rect 4291 429 4293 433
rect 4297 429 4299 433
rect 4303 429 4305 433
rect 4309 429 4311 433
rect 4315 429 4317 433
rect 4321 429 4323 433
rect 4327 429 4465 433
rect 4469 429 4471 433
rect 4475 429 4477 433
rect 4481 429 4483 433
rect 4487 429 4489 433
rect 4493 429 4495 433
rect 4499 429 4501 433
rect 4505 429 4589 433
rect 411 427 4589 429
rect 411 423 495 427
rect 499 423 501 427
rect 505 423 507 427
rect 511 423 513 427
rect 517 423 519 427
rect 523 423 525 427
rect 529 423 531 427
rect 535 423 673 427
rect 677 423 679 427
rect 683 423 685 427
rect 689 423 691 427
rect 695 423 697 427
rect 701 423 703 427
rect 707 423 709 427
rect 713 423 969 427
rect 973 423 975 427
rect 979 423 981 427
rect 985 423 987 427
rect 991 423 993 427
rect 997 423 999 427
rect 1003 423 1005 427
rect 1009 423 1147 427
rect 1151 423 1153 427
rect 1157 423 1159 427
rect 1163 423 1165 427
rect 1169 423 1171 427
rect 1175 423 1177 427
rect 1181 423 1183 427
rect 1187 423 1443 427
rect 1447 423 1449 427
rect 1453 423 1455 427
rect 1459 423 1461 427
rect 1465 423 1467 427
rect 1471 423 1473 427
rect 1477 423 1479 427
rect 1483 423 1621 427
rect 1625 423 1627 427
rect 1631 423 1633 427
rect 1637 423 1639 427
rect 1643 423 1645 427
rect 1649 423 1651 427
rect 1655 423 1657 427
rect 1661 423 1917 427
rect 1921 423 1923 427
rect 1927 423 1929 427
rect 1933 423 1935 427
rect 1939 423 1941 427
rect 1945 423 1947 427
rect 1951 423 1953 427
rect 1957 423 2095 427
rect 2099 423 2101 427
rect 2105 423 2107 427
rect 2111 423 2113 427
rect 2117 423 2119 427
rect 2123 423 2125 427
rect 2129 423 2131 427
rect 2135 423 2391 427
rect 2395 423 2397 427
rect 2401 423 2403 427
rect 2407 423 2409 427
rect 2413 423 2415 427
rect 2419 423 2421 427
rect 2425 423 2427 427
rect 2431 423 2569 427
rect 2573 423 2575 427
rect 2579 423 2581 427
rect 2585 423 2587 427
rect 2591 423 2593 427
rect 2597 423 2599 427
rect 2603 423 2605 427
rect 2609 423 2865 427
rect 2869 423 2871 427
rect 2875 423 2877 427
rect 2881 423 2883 427
rect 2887 423 2889 427
rect 2893 423 2895 427
rect 2899 423 2901 427
rect 2905 423 3043 427
rect 3047 423 3049 427
rect 3053 423 3055 427
rect 3059 423 3061 427
rect 3065 423 3067 427
rect 3071 423 3073 427
rect 3077 423 3079 427
rect 3083 423 3339 427
rect 3343 423 3345 427
rect 3349 423 3351 427
rect 3355 423 3357 427
rect 3361 423 3363 427
rect 3367 423 3369 427
rect 3373 423 3375 427
rect 3379 423 3517 427
rect 3521 423 3523 427
rect 3527 423 3529 427
rect 3533 423 3535 427
rect 3539 423 3541 427
rect 3545 423 3547 427
rect 3551 423 3553 427
rect 3557 423 3813 427
rect 3817 423 3819 427
rect 3823 423 3825 427
rect 3829 423 3831 427
rect 3835 423 3837 427
rect 3841 423 3843 427
rect 3847 423 3849 427
rect 3853 423 3991 427
rect 3995 423 3997 427
rect 4001 423 4003 427
rect 4007 423 4009 427
rect 4013 423 4015 427
rect 4019 423 4021 427
rect 4025 423 4027 427
rect 4031 423 4287 427
rect 4291 423 4293 427
rect 4297 423 4299 427
rect 4303 423 4305 427
rect 4309 423 4311 427
rect 4315 423 4317 427
rect 4321 423 4323 427
rect 4327 423 4465 427
rect 4469 423 4471 427
rect 4475 423 4477 427
rect 4481 423 4483 427
rect 4487 423 4489 427
rect 4493 423 4495 427
rect 4499 423 4501 427
rect 4505 423 4589 427
rect 411 421 4589 423
rect 411 412 495 421
rect 499 412 501 421
rect 505 412 507 421
rect 511 412 513 421
rect 517 412 519 421
rect 523 412 525 421
rect 529 412 531 421
rect 535 412 673 421
rect 677 412 679 421
rect 683 412 685 421
rect 689 412 691 421
rect 695 412 697 421
rect 701 412 703 421
rect 707 412 709 421
rect 713 412 969 421
rect 973 412 975 421
rect 979 412 981 421
rect 985 412 987 421
rect 991 412 993 421
rect 997 412 999 421
rect 1003 412 1005 421
rect 1009 412 1147 421
rect 1151 412 1153 421
rect 1157 412 1159 421
rect 1163 412 1165 421
rect 1169 412 1171 421
rect 1175 412 1177 421
rect 1181 412 1183 421
rect 1187 412 1443 421
rect 1447 412 1449 421
rect 1453 412 1455 421
rect 1459 412 1461 421
rect 1465 412 1467 421
rect 1471 412 1473 421
rect 1477 412 1479 421
rect 1483 412 1621 421
rect 1625 412 1627 421
rect 1631 412 1633 421
rect 1637 412 1639 421
rect 1643 412 1645 421
rect 1649 412 1651 421
rect 1655 412 1657 421
rect 1661 412 1917 421
rect 1921 412 1923 421
rect 1927 412 1929 421
rect 1933 412 1935 421
rect 1939 412 1941 421
rect 1945 412 1947 421
rect 1951 412 1953 421
rect 1957 412 2095 421
rect 2099 412 2101 421
rect 2105 412 2107 421
rect 2111 412 2113 421
rect 2117 412 2119 421
rect 2123 412 2125 421
rect 2129 412 2131 421
rect 2135 412 2391 421
rect 2395 412 2397 421
rect 2401 412 2403 421
rect 2407 412 2409 421
rect 2413 412 2415 421
rect 2419 412 2421 421
rect 2425 412 2427 421
rect 2431 412 2569 421
rect 2573 412 2575 421
rect 2579 412 2581 421
rect 2585 412 2587 421
rect 2591 412 2593 421
rect 2597 412 2599 421
rect 2603 412 2605 421
rect 2609 412 2865 421
rect 2869 412 2871 421
rect 2875 412 2877 421
rect 2881 412 2883 421
rect 2887 412 2889 421
rect 2893 412 2895 421
rect 2899 412 2901 421
rect 2905 412 3043 421
rect 3047 412 3049 421
rect 3053 412 3055 421
rect 3059 412 3061 421
rect 3065 412 3067 421
rect 3071 412 3073 421
rect 3077 412 3079 421
rect 3083 412 3339 421
rect 3343 412 3345 421
rect 3349 412 3351 421
rect 3355 412 3357 421
rect 3361 412 3363 421
rect 3367 412 3369 421
rect 3373 412 3375 421
rect 3379 412 3517 421
rect 3521 412 3523 421
rect 3527 412 3529 421
rect 3533 412 3535 421
rect 3539 412 3541 421
rect 3545 412 3547 421
rect 3551 412 3553 421
rect 3557 412 3813 421
rect 3817 412 3819 421
rect 3823 412 3825 421
rect 3829 412 3831 421
rect 3835 412 3837 421
rect 3841 412 3843 421
rect 3847 412 3849 421
rect 3853 412 3991 421
rect 3995 412 3997 421
rect 4001 412 4003 421
rect 4007 412 4009 421
rect 4013 412 4015 421
rect 4019 412 4021 421
rect 4025 412 4027 421
rect 4031 412 4287 421
rect 4291 412 4293 421
rect 4297 412 4299 421
rect 4303 412 4305 421
rect 4309 412 4311 421
rect 4315 412 4317 421
rect 4321 412 4323 421
rect 4327 412 4465 421
rect 4469 412 4471 421
rect 4475 412 4477 421
rect 4481 412 4483 421
rect 4487 412 4489 421
rect 4493 412 4495 421
rect 4499 412 4501 421
rect 4505 412 4589 421
rect 411 411 4589 412
rect 367 406 4633 407
rect 367 402 539 406
rect 543 402 545 406
rect 549 402 551 406
rect 555 402 557 406
rect 561 402 563 406
rect 567 402 569 406
rect 573 402 575 406
rect 579 402 629 406
rect 633 402 635 406
rect 639 402 641 406
rect 645 402 647 406
rect 651 402 653 406
rect 657 402 659 406
rect 663 402 665 406
rect 669 402 1013 406
rect 1017 402 1019 406
rect 1023 402 1025 406
rect 1029 402 1031 406
rect 1035 402 1037 406
rect 1041 402 1043 406
rect 1047 402 1049 406
rect 1053 402 1103 406
rect 1107 402 1109 406
rect 1113 402 1115 406
rect 1119 402 1121 406
rect 1125 402 1127 406
rect 1131 402 1133 406
rect 1137 402 1139 406
rect 1143 402 1487 406
rect 1491 402 1493 406
rect 1497 402 1499 406
rect 1503 402 1505 406
rect 1509 402 1511 406
rect 1515 402 1517 406
rect 1521 402 1523 406
rect 1527 402 1577 406
rect 1581 402 1583 406
rect 1587 402 1589 406
rect 1593 402 1595 406
rect 1599 402 1601 406
rect 1605 402 1607 406
rect 1611 402 1613 406
rect 1617 402 1961 406
rect 1965 402 1967 406
rect 1971 402 1973 406
rect 1977 402 1979 406
rect 1983 402 1985 406
rect 1989 402 1991 406
rect 1995 402 1997 406
rect 2001 402 2051 406
rect 2055 402 2057 406
rect 2061 402 2063 406
rect 2067 402 2069 406
rect 2073 402 2075 406
rect 2079 402 2081 406
rect 2085 402 2087 406
rect 2091 402 2435 406
rect 2439 402 2441 406
rect 2445 402 2447 406
rect 2451 402 2453 406
rect 2457 402 2459 406
rect 2463 402 2465 406
rect 2469 402 2471 406
rect 2475 402 2525 406
rect 2529 402 2531 406
rect 2535 402 2537 406
rect 2541 402 2543 406
rect 2547 402 2549 406
rect 2553 402 2555 406
rect 2559 402 2561 406
rect 2565 402 2909 406
rect 2913 402 2915 406
rect 2919 402 2921 406
rect 2925 402 2927 406
rect 2931 402 2933 406
rect 2937 402 2939 406
rect 2943 402 2945 406
rect 2949 402 2999 406
rect 3003 402 3005 406
rect 3009 402 3011 406
rect 3015 402 3017 406
rect 3021 402 3023 406
rect 3027 402 3029 406
rect 3033 402 3035 406
rect 3039 402 3383 406
rect 3387 402 3389 406
rect 3393 402 3395 406
rect 3399 402 3401 406
rect 3405 402 3407 406
rect 3411 402 3413 406
rect 3417 402 3419 406
rect 3423 402 3473 406
rect 3477 402 3479 406
rect 3483 402 3485 406
rect 3489 402 3491 406
rect 3495 402 3497 406
rect 3501 402 3503 406
rect 3507 402 3509 406
rect 3513 402 3857 406
rect 3861 402 3863 406
rect 3867 402 3869 406
rect 3873 402 3875 406
rect 3879 402 3881 406
rect 3885 402 3887 406
rect 3891 402 3893 406
rect 3897 402 3947 406
rect 3951 402 3953 406
rect 3957 402 3959 406
rect 3963 402 3965 406
rect 3969 402 3971 406
rect 3975 402 3977 406
rect 3981 402 3983 406
rect 3987 402 4331 406
rect 4335 402 4337 406
rect 4341 402 4343 406
rect 4347 402 4349 406
rect 4353 402 4355 406
rect 4359 402 4361 406
rect 4365 402 4367 406
rect 4371 402 4421 406
rect 4425 402 4427 406
rect 4431 402 4433 406
rect 4437 402 4439 406
rect 4443 402 4445 406
rect 4449 402 4451 406
rect 4455 402 4457 406
rect 4461 402 4516 406
rect 4520 402 4522 406
rect 4526 402 4528 406
rect 4532 402 4534 406
rect 4538 402 4540 406
rect 4544 402 4546 406
rect 4550 402 4552 406
rect 4556 402 4558 406
rect 4562 402 4564 406
rect 4568 402 4570 406
rect 4574 402 4576 406
rect 4580 402 4582 406
rect 4586 402 4588 406
rect 4592 402 4594 406
rect 4598 402 4600 406
rect 4604 402 4606 406
rect 4610 402 4612 406
rect 4616 402 4618 406
rect 4622 402 4633 406
rect 367 400 4633 402
rect 367 396 4516 400
rect 4520 396 4522 400
rect 4526 396 4528 400
rect 4532 396 4534 400
rect 4538 396 4540 400
rect 4544 396 4546 400
rect 4550 396 4552 400
rect 4556 396 4558 400
rect 4562 396 4564 400
rect 4568 396 4570 400
rect 4574 396 4576 400
rect 4580 396 4582 400
rect 4586 396 4588 400
rect 4592 396 4594 400
rect 4598 396 4600 400
rect 4604 396 4606 400
rect 4610 396 4612 400
rect 4616 396 4618 400
rect 4622 396 4633 400
rect 367 394 4633 396
rect 367 390 539 394
rect 543 390 545 394
rect 549 390 551 394
rect 555 390 557 394
rect 561 390 563 394
rect 567 390 569 394
rect 573 390 575 394
rect 579 390 629 394
rect 633 390 635 394
rect 639 390 641 394
rect 645 390 647 394
rect 651 390 653 394
rect 657 390 659 394
rect 663 390 665 394
rect 669 390 1013 394
rect 1017 390 1019 394
rect 1023 390 1025 394
rect 1029 390 1031 394
rect 1035 390 1037 394
rect 1041 390 1043 394
rect 1047 390 1049 394
rect 1053 390 1103 394
rect 1107 390 1109 394
rect 1113 390 1115 394
rect 1119 390 1121 394
rect 1125 390 1127 394
rect 1131 390 1133 394
rect 1137 390 1139 394
rect 1143 390 1487 394
rect 1491 390 1493 394
rect 1497 390 1499 394
rect 1503 390 1505 394
rect 1509 390 1511 394
rect 1515 390 1517 394
rect 1521 390 1523 394
rect 1527 390 1577 394
rect 1581 390 1583 394
rect 1587 390 1589 394
rect 1593 390 1595 394
rect 1599 390 1601 394
rect 1605 390 1607 394
rect 1611 390 1613 394
rect 1617 390 1961 394
rect 1965 390 1967 394
rect 1971 390 1973 394
rect 1977 390 1979 394
rect 1983 390 1985 394
rect 1989 390 1991 394
rect 1995 390 1997 394
rect 2001 390 2051 394
rect 2055 390 2057 394
rect 2061 390 2063 394
rect 2067 390 2069 394
rect 2073 390 2075 394
rect 2079 390 2081 394
rect 2085 390 2087 394
rect 2091 390 2435 394
rect 2439 390 2441 394
rect 2445 390 2447 394
rect 2451 390 2453 394
rect 2457 390 2459 394
rect 2463 390 2465 394
rect 2469 390 2471 394
rect 2475 390 2525 394
rect 2529 390 2531 394
rect 2535 390 2537 394
rect 2541 390 2543 394
rect 2547 390 2549 394
rect 2553 390 2555 394
rect 2559 390 2561 394
rect 2565 390 2909 394
rect 2913 390 2915 394
rect 2919 390 2921 394
rect 2925 390 2927 394
rect 2931 390 2933 394
rect 2937 390 2939 394
rect 2943 390 2945 394
rect 2949 390 2999 394
rect 3003 390 3005 394
rect 3009 390 3011 394
rect 3015 390 3017 394
rect 3021 390 3023 394
rect 3027 390 3029 394
rect 3033 390 3035 394
rect 3039 390 3383 394
rect 3387 390 3389 394
rect 3393 390 3395 394
rect 3399 390 3401 394
rect 3405 390 3407 394
rect 3411 390 3413 394
rect 3417 390 3419 394
rect 3423 390 3473 394
rect 3477 390 3479 394
rect 3483 390 3485 394
rect 3489 390 3491 394
rect 3495 390 3497 394
rect 3501 390 3503 394
rect 3507 390 3509 394
rect 3513 390 3857 394
rect 3861 390 3863 394
rect 3867 390 3869 394
rect 3873 390 3875 394
rect 3879 390 3881 394
rect 3885 390 3887 394
rect 3891 390 3893 394
rect 3897 390 3947 394
rect 3951 390 3953 394
rect 3957 390 3959 394
rect 3963 390 3965 394
rect 3969 390 3971 394
rect 3975 390 3977 394
rect 3981 390 3983 394
rect 3987 390 4331 394
rect 4335 390 4337 394
rect 4341 390 4343 394
rect 4347 390 4349 394
rect 4353 390 4355 394
rect 4359 390 4361 394
rect 4365 390 4367 394
rect 4371 390 4421 394
rect 4425 390 4427 394
rect 4431 390 4433 394
rect 4437 390 4439 394
rect 4443 390 4445 394
rect 4449 390 4451 394
rect 4455 390 4457 394
rect 4461 390 4516 394
rect 4520 390 4522 394
rect 4526 390 4528 394
rect 4532 390 4534 394
rect 4538 390 4540 394
rect 4544 390 4546 394
rect 4550 390 4552 394
rect 4556 390 4558 394
rect 4562 390 4564 394
rect 4568 390 4570 394
rect 4574 390 4576 394
rect 4580 390 4582 394
rect 4586 390 4588 394
rect 4592 390 4594 394
rect 4598 390 4600 394
rect 4604 390 4606 394
rect 4610 390 4612 394
rect 4616 390 4618 394
rect 4622 390 4633 394
rect 367 388 4633 390
rect 367 384 4516 388
rect 4520 384 4522 388
rect 4526 384 4528 388
rect 4532 384 4534 388
rect 4538 384 4540 388
rect 4544 384 4546 388
rect 4550 384 4552 388
rect 4556 384 4558 388
rect 4562 384 4564 388
rect 4568 384 4570 388
rect 4574 384 4576 388
rect 4580 384 4582 388
rect 4586 384 4588 388
rect 4592 384 4594 388
rect 4598 384 4600 388
rect 4604 384 4606 388
rect 4610 384 4612 388
rect 4616 384 4618 388
rect 4622 384 4633 388
rect 367 382 4633 384
rect 367 378 545 382
rect 549 378 551 382
rect 555 378 557 382
rect 561 378 563 382
rect 567 378 569 382
rect 573 378 575 382
rect 579 378 629 382
rect 633 378 635 382
rect 639 378 641 382
rect 645 378 647 382
rect 651 378 653 382
rect 657 378 659 382
rect 663 378 1019 382
rect 1023 378 1025 382
rect 1029 378 1031 382
rect 1035 378 1037 382
rect 1041 378 1043 382
rect 1047 378 1049 382
rect 1053 378 1103 382
rect 1107 378 1109 382
rect 1113 378 1115 382
rect 1119 378 1121 382
rect 1125 378 1127 382
rect 1131 378 1133 382
rect 1137 378 1493 382
rect 1497 378 1499 382
rect 1503 378 1505 382
rect 1509 378 1511 382
rect 1515 378 1517 382
rect 1521 378 1523 382
rect 1527 378 1577 382
rect 1581 378 1583 382
rect 1587 378 1589 382
rect 1593 378 1595 382
rect 1599 378 1601 382
rect 1605 378 1607 382
rect 1611 378 1967 382
rect 1971 378 1973 382
rect 1977 378 1979 382
rect 1983 378 1985 382
rect 1989 378 1991 382
rect 1995 378 1997 382
rect 2001 378 2051 382
rect 2055 378 2057 382
rect 2061 378 2063 382
rect 2067 378 2069 382
rect 2073 378 2075 382
rect 2079 378 2081 382
rect 2085 378 2441 382
rect 2445 378 2447 382
rect 2451 378 2453 382
rect 2457 378 2459 382
rect 2463 378 2465 382
rect 2469 378 2471 382
rect 2475 378 2525 382
rect 2529 378 2531 382
rect 2535 378 2537 382
rect 2541 378 2543 382
rect 2547 378 2549 382
rect 2553 378 2555 382
rect 2559 378 2915 382
rect 2919 378 2921 382
rect 2925 378 2927 382
rect 2931 378 2933 382
rect 2937 378 2939 382
rect 2943 378 2945 382
rect 2949 378 2999 382
rect 3003 378 3005 382
rect 3009 378 3011 382
rect 3015 378 3017 382
rect 3021 378 3023 382
rect 3027 378 3029 382
rect 3033 378 3389 382
rect 3393 378 3395 382
rect 3399 378 3401 382
rect 3405 378 3407 382
rect 3411 378 3413 382
rect 3417 378 3419 382
rect 3423 378 3473 382
rect 3477 378 3479 382
rect 3483 378 3485 382
rect 3489 378 3491 382
rect 3495 378 3497 382
rect 3501 378 3503 382
rect 3507 378 3863 382
rect 3867 378 3869 382
rect 3873 378 3875 382
rect 3879 378 3881 382
rect 3885 378 3887 382
rect 3891 378 3893 382
rect 3897 378 3947 382
rect 3951 378 3953 382
rect 3957 378 3959 382
rect 3963 378 3965 382
rect 3969 378 3971 382
rect 3975 378 3977 382
rect 3981 378 4337 382
rect 4341 378 4343 382
rect 4347 378 4349 382
rect 4353 378 4355 382
rect 4359 378 4361 382
rect 4365 378 4367 382
rect 4371 378 4421 382
rect 4425 378 4427 382
rect 4431 378 4433 382
rect 4437 378 4439 382
rect 4443 378 4445 382
rect 4449 378 4451 382
rect 4455 378 4516 382
rect 4520 378 4522 382
rect 4526 378 4528 382
rect 4532 378 4534 382
rect 4538 378 4540 382
rect 4544 378 4546 382
rect 4550 378 4552 382
rect 4556 378 4558 382
rect 4562 378 4564 382
rect 4568 378 4570 382
rect 4574 378 4576 382
rect 4580 378 4582 382
rect 4586 378 4588 382
rect 4592 378 4594 382
rect 4598 378 4600 382
rect 4604 378 4606 382
rect 4610 378 4612 382
rect 4616 378 4618 382
rect 4622 378 4633 382
rect 367 367 4633 378
rect 320 259 356 260
rect 320 255 321 259
rect 325 255 327 259
rect 331 255 333 259
rect 337 255 339 259
rect 343 255 345 259
rect 349 255 351 259
rect 355 255 356 259
rect 320 247 356 255
rect 320 243 321 247
rect 325 243 327 247
rect 331 243 333 247
rect 337 243 339 247
rect 343 243 345 247
rect 349 243 351 247
rect 355 243 356 247
rect 320 235 356 243
rect 320 231 321 235
rect 325 231 327 235
rect 331 231 333 235
rect 337 231 339 235
rect 343 231 345 235
rect 349 231 351 235
rect 355 231 356 235
rect 320 223 356 231
rect 320 219 321 223
rect 325 219 327 223
rect 331 219 333 223
rect 337 219 339 223
rect 343 219 345 223
rect 349 219 351 223
rect 355 219 356 223
rect 320 218 356 219
rect 4644 259 4680 260
rect 4644 255 4645 259
rect 4649 255 4651 259
rect 4655 255 4657 259
rect 4661 255 4663 259
rect 4667 255 4669 259
rect 4673 255 4675 259
rect 4679 255 4680 259
rect 4644 247 4680 255
rect 4644 243 4645 247
rect 4649 243 4651 247
rect 4655 243 4657 247
rect 4661 243 4663 247
rect 4667 243 4669 247
rect 4673 243 4675 247
rect 4679 243 4680 247
rect 4644 235 4680 243
rect 4644 231 4645 235
rect 4649 231 4651 235
rect 4655 231 4657 235
rect 4661 231 4663 235
rect 4667 231 4669 235
rect 4673 231 4675 235
rect 4679 231 4680 235
rect 4644 223 4680 231
rect 4644 219 4645 223
rect 4649 219 4651 223
rect 4655 219 4657 223
rect 4661 219 4663 223
rect 4667 219 4669 223
rect 4673 219 4675 223
rect 4679 219 4680 223
rect 4644 218 4680 219
<< m3contact >>
rect 467 467 531 496
rect 4516 402 4520 406
rect 4522 402 4526 406
rect 4528 402 4532 406
rect 4534 402 4538 406
rect 4540 402 4544 406
rect 4546 402 4550 406
rect 4552 402 4556 406
rect 4558 402 4562 406
rect 4564 402 4568 406
rect 4570 402 4574 406
rect 4576 402 4580 406
rect 4582 402 4586 406
rect 4588 402 4592 406
rect 4594 402 4598 406
rect 4600 402 4604 406
rect 4606 402 4610 406
rect 4612 402 4616 406
rect 4618 402 4622 406
rect 4516 396 4520 400
rect 4522 396 4526 400
rect 4528 396 4532 400
rect 4534 396 4538 400
rect 4540 396 4544 400
rect 4546 396 4550 400
rect 4552 396 4556 400
rect 4558 396 4562 400
rect 4564 396 4568 400
rect 4570 396 4574 400
rect 4576 396 4580 400
rect 4582 396 4586 400
rect 4588 396 4592 400
rect 4594 396 4598 400
rect 4600 396 4604 400
rect 4606 396 4610 400
rect 4612 396 4616 400
rect 4618 396 4622 400
rect 4516 390 4520 394
rect 4522 390 4526 394
rect 4528 390 4532 394
rect 4534 390 4538 394
rect 4540 390 4544 394
rect 4546 390 4550 394
rect 4552 390 4556 394
rect 4558 390 4562 394
rect 4564 390 4568 394
rect 4570 390 4574 394
rect 4576 390 4580 394
rect 4582 390 4586 394
rect 4588 390 4592 394
rect 4594 390 4598 394
rect 4600 390 4604 394
rect 4606 390 4610 394
rect 4612 390 4616 394
rect 4618 390 4622 394
rect 4516 384 4520 388
rect 4522 384 4526 388
rect 4528 384 4532 388
rect 4534 384 4538 388
rect 4540 384 4544 388
rect 4546 384 4550 388
rect 4552 384 4556 388
rect 4558 384 4562 388
rect 4564 384 4568 388
rect 4570 384 4574 388
rect 4576 384 4580 388
rect 4582 384 4586 388
rect 4588 384 4592 388
rect 4594 384 4598 388
rect 4600 384 4604 388
rect 4606 384 4610 388
rect 4612 384 4616 388
rect 4618 384 4622 388
rect 4516 378 4520 382
rect 4522 378 4526 382
rect 4528 378 4532 382
rect 4534 378 4538 382
rect 4540 378 4544 382
rect 4546 378 4550 382
rect 4552 378 4556 382
rect 4558 378 4562 382
rect 4564 378 4568 382
rect 4570 378 4574 382
rect 4576 378 4580 382
rect 4582 378 4586 382
rect 4588 378 4592 382
rect 4594 378 4598 382
rect 4600 378 4604 382
rect 4606 378 4610 382
rect 4612 378 4616 382
rect 4618 378 4622 382
rect 321 255 325 259
rect 333 255 337 259
rect 345 255 349 259
rect 327 243 331 247
rect 339 243 343 247
rect 351 243 355 247
rect 321 231 325 235
rect 333 231 337 235
rect 345 231 349 235
rect 327 219 331 223
rect 339 219 343 223
rect 351 219 355 223
rect 4651 255 4655 259
rect 4663 255 4667 259
rect 4675 255 4679 259
rect 4645 243 4649 247
rect 4657 243 4661 247
rect 4669 243 4673 247
rect 4651 231 4655 235
rect 4663 231 4667 235
rect 4675 231 4679 235
rect 4645 219 4649 223
rect 4657 219 4661 223
rect 4669 219 4673 223
<< metal3 >>
rect 347 496 532 497
rect 347 467 467 496
rect 531 467 532 496
rect 347 466 532 467
rect 347 260 387 466
rect 4515 406 4653 407
rect 4515 402 4516 406
rect 4520 402 4522 406
rect 4526 402 4528 406
rect 4532 402 4534 406
rect 4538 402 4540 406
rect 4544 402 4546 406
rect 4550 402 4552 406
rect 4556 402 4558 406
rect 4562 402 4564 406
rect 4568 402 4570 406
rect 4574 402 4576 406
rect 4580 402 4582 406
rect 4586 402 4588 406
rect 4592 402 4594 406
rect 4598 402 4600 406
rect 4604 402 4606 406
rect 4610 402 4612 406
rect 4616 402 4618 406
rect 4622 402 4653 406
rect 4515 400 4653 402
rect 4515 396 4516 400
rect 4520 396 4522 400
rect 4526 396 4528 400
rect 4532 396 4534 400
rect 4538 396 4540 400
rect 4544 396 4546 400
rect 4550 396 4552 400
rect 4556 396 4558 400
rect 4562 396 4564 400
rect 4568 396 4570 400
rect 4574 396 4576 400
rect 4580 396 4582 400
rect 4586 396 4588 400
rect 4592 396 4594 400
rect 4598 396 4600 400
rect 4604 396 4606 400
rect 4610 396 4612 400
rect 4616 396 4618 400
rect 4622 396 4653 400
rect 4515 394 4653 396
rect 4515 390 4516 394
rect 4520 390 4522 394
rect 4526 390 4528 394
rect 4532 390 4534 394
rect 4538 390 4540 394
rect 4544 390 4546 394
rect 4550 390 4552 394
rect 4556 390 4558 394
rect 4562 390 4564 394
rect 4568 390 4570 394
rect 4574 390 4576 394
rect 4580 390 4582 394
rect 4586 390 4588 394
rect 4592 390 4594 394
rect 4598 390 4600 394
rect 4604 390 4606 394
rect 4610 390 4612 394
rect 4616 390 4618 394
rect 4622 390 4653 394
rect 4515 388 4653 390
rect 4515 384 4516 388
rect 4520 384 4522 388
rect 4526 384 4528 388
rect 4532 384 4534 388
rect 4538 384 4540 388
rect 4544 384 4546 388
rect 4550 384 4552 388
rect 4556 384 4558 388
rect 4562 384 4564 388
rect 4568 384 4570 388
rect 4574 384 4576 388
rect 4580 384 4582 388
rect 4586 384 4588 388
rect 4592 384 4594 388
rect 4598 384 4600 388
rect 4604 384 4606 388
rect 4610 384 4612 388
rect 4616 384 4618 388
rect 4622 384 4653 388
rect 4515 382 4653 384
rect 4515 378 4516 382
rect 4520 378 4522 382
rect 4526 378 4528 382
rect 4532 378 4534 382
rect 4538 378 4540 382
rect 4544 378 4546 382
rect 4550 378 4552 382
rect 4556 378 4558 382
rect 4562 378 4564 382
rect 4568 378 4570 382
rect 4574 378 4576 382
rect 4580 378 4582 382
rect 4586 378 4588 382
rect 4592 378 4594 382
rect 4598 378 4600 382
rect 4604 378 4606 382
rect 4610 378 4612 382
rect 4616 378 4618 382
rect 4622 378 4653 382
rect 4515 376 4653 378
rect 260 259 387 260
rect 260 255 321 259
rect 325 255 333 259
rect 337 255 345 259
rect 349 255 387 259
rect 260 247 387 255
rect 260 243 327 247
rect 331 243 339 247
rect 343 243 351 247
rect 355 243 387 247
rect 260 235 387 243
rect 260 231 321 235
rect 325 231 333 235
rect 337 231 345 235
rect 349 231 387 235
rect 260 223 387 231
rect 260 219 327 223
rect 331 219 339 223
rect 343 219 351 223
rect 355 219 387 223
rect 260 0 387 219
rect 4613 260 4653 376
rect 4613 259 4740 260
rect 4613 255 4651 259
rect 4655 255 4663 259
rect 4667 255 4675 259
rect 4679 255 4740 259
rect 4613 247 4740 255
rect 4613 243 4645 247
rect 4649 243 4657 247
rect 4661 243 4669 247
rect 4673 243 4740 247
rect 4613 235 4740 243
rect 4613 231 4651 235
rect 4655 231 4663 235
rect 4667 231 4675 235
rect 4679 231 4740 235
rect 4613 223 4740 231
rect 4613 219 4645 223
rect 4649 219 4657 223
rect 4661 219 4669 223
rect 4673 219 4740 223
rect 4613 0 4740 219
use bondingpad  bondingpad_1
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 260 260
use bondingpad  bondingpad_0
timestamp 1259953556
transform 1 0 4740 0 1 0
box 0 0 260 260
<< labels >>
rlabel m2contact 4307 512 4307 512 6 Gnd
rlabel m2contact 4441 512 4441 512 6 CVdd
rlabel m2contact 4412 512 4412 512 6 Bias
rlabel m2contact 4379 512 4379 512 6 Bias
rlabel m2contact 4351 512 4351 512 6 CVdd
rlabel m2contact 3833 512 3833 512 6 Gnd
rlabel m2contact 4011 512 4011 512 6 Gnd
rlabel m2contact 3967 512 3967 512 6 CVdd
rlabel m2contact 3938 512 3938 512 6 Bias
rlabel m2contact 3905 512 3905 512 6 Bias
rlabel m2contact 3877 512 3877 512 6 CVdd
rlabel m2contact 3359 512 3359 512 6 Gnd
rlabel m2contact 3537 512 3537 512 6 Gnd
rlabel m2contact 3493 512 3493 512 6 CVdd
rlabel m2contact 3464 512 3464 512 6 Bias
rlabel m2contact 3431 512 3431 512 6 Bias
rlabel m2contact 3403 512 3403 512 6 CVdd
rlabel m2contact 2885 512 2885 512 6 Gnd
rlabel m2contact 3063 512 3063 512 6 Gnd
rlabel m2contact 3019 512 3019 512 6 CVdd
rlabel m2contact 2990 512 2990 512 6 Bias
rlabel m2contact 2957 512 2957 512 6 Bias
rlabel m2contact 2929 512 2929 512 6 CVdd
rlabel m2contact 2411 512 2411 512 6 Gnd
rlabel m2contact 2589 512 2589 512 6 Gnd
rlabel m2contact 2545 512 2545 512 6 CVdd
rlabel m2contact 2516 512 2516 512 6 Bias
rlabel m2contact 2483 512 2483 512 6 Bias
rlabel m2contact 2455 512 2455 512 6 CVdd
rlabel m2contact 1937 512 1937 512 6 Gnd
rlabel m2contact 2115 512 2115 512 6 Gnd
rlabel m2contact 2071 512 2071 512 6 CVdd
rlabel m2contact 2042 512 2042 512 6 Bias
rlabel m2contact 2009 512 2009 512 6 Bias
rlabel m2contact 1981 512 1981 512 6 CVdd
rlabel m2contact 1463 512 1463 512 6 Gnd
rlabel m2contact 1641 512 1641 512 6 Gnd
rlabel m2contact 1597 512 1597 512 6 CVdd
rlabel m2contact 1568 512 1568 512 6 Bias
rlabel m2contact 1535 512 1535 512 6 Bias
rlabel m2contact 1507 512 1507 512 6 CVdd
rlabel m2contact 989 512 989 512 6 Gnd
rlabel m2contact 1167 512 1167 512 6 Gnd
rlabel m2contact 1123 512 1123 512 6 CVdd
rlabel m2contact 1094 512 1094 512 6 Bias
rlabel m2contact 1061 512 1061 512 6 Bias
rlabel m2contact 1033 512 1033 512 6 CVdd
rlabel m2contact 693 512 693 512 6 Gnd
rlabel m2contact 649 512 649 512 6 CVdd
rlabel m2contact 620 512 620 512 6 Bias
rlabel m2contact 587 512 587 512 6 Bias
rlabel m2contact 559 512 559 512 6 CVdd
<< end >>
