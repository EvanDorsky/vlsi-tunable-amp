magic
tech scmos
timestamp 1418846892
<< ntransistor >>
rect -5 -138 -1 -136
rect 6 -138 10 -136
rect 0 -145 4 -143
rect 2 -168 4 -164
<< ptransistor >>
rect -5 -88 -1 -86
rect 6 -88 10 -86
rect -5 -108 -1 -106
rect 6 -108 10 -106
rect 2 -184 4 -180
<< ndiffusion >>
rect -5 -136 -1 -135
rect 6 -136 10 -135
rect -5 -139 -1 -138
rect 6 -139 10 -138
rect -5 -142 10 -139
rect 0 -143 4 -142
rect 0 -146 4 -145
rect -1 -149 6 -146
rect 1 -168 2 -164
rect 4 -168 5 -164
<< pdiffusion >>
rect -5 -86 -1 -85
rect 6 -86 10 -85
rect -5 -89 -1 -88
rect 6 -89 10 -88
rect -5 -106 -1 -105
rect 6 -106 10 -105
rect -5 -109 -1 -108
rect 6 -109 10 -108
rect 1 -184 2 -180
rect 4 -184 5 -180
<< ndcontact >>
rect -5 -135 -1 -131
rect 6 -135 10 -131
rect -5 -150 -1 -146
rect 6 -150 10 -146
rect -3 -168 1 -164
rect 5 -168 9 -164
<< pdcontact >>
rect -5 -85 -1 -81
rect 6 -85 10 -81
rect -5 -93 -1 -89
rect 6 -93 10 -89
rect -5 -105 -1 -101
rect 6 -105 10 -101
rect -5 -113 -1 -109
rect 6 -113 10 -109
rect -3 -184 1 -180
rect 5 -184 9 -180
<< polysilicon >>
rect -10 -88 -5 -86
rect -1 -88 6 -86
rect 10 -88 14 -86
rect -8 -108 -5 -106
rect -1 -108 1 -106
rect 4 -108 6 -106
rect 10 -108 13 -106
rect -8 -126 -6 -108
rect 11 -116 13 -108
rect 3 -118 13 -116
rect -8 -128 2 -126
rect -8 -136 -6 -128
rect 11 -136 13 -118
rect -8 -138 -5 -136
rect -1 -138 1 -136
rect 4 -138 6 -136
rect 10 -138 13 -136
rect -10 -145 0 -143
rect 4 -145 14 -143
rect 2 -164 4 -161
rect 2 -180 4 -168
rect 2 -186 4 -184
<< polycontact >>
rect -1 -119 3 -115
rect 2 -129 6 -125
rect 2 -161 6 -157
<< metal1 >>
rect -5 -94 -1 -93
rect 6 -94 10 -93
rect -10 -105 -5 -101
rect -1 -105 6 -101
rect 10 -105 14 -101
rect -5 -120 -1 -113
rect -5 -131 -1 -124
rect 6 -120 10 -113
rect 6 -131 10 -124
rect -10 -146 14 -145
rect -10 -149 -5 -146
rect -1 -149 6 -146
rect 10 -149 14 -146
rect -3 -180 1 -168
<< m2contact >>
rect -5 -98 -1 -94
rect 6 -98 10 -94
rect -5 -124 -1 -120
rect 6 -124 10 -120
rect 2 -157 6 -153
<< metal2 >>
rect -5 -120 -1 -98
rect 6 -120 10 -98
rect 2 -153 6 -120
<< labels >>
rlabel metal1 13 -149 14 -145 8 Gnd
rlabel metal1 -10 -105 -9 -101 3 Vdd
rlabel m2contact 6 -98 10 -94 1 Qbar
rlabel pdcontact 6 -85 10 -81 1 Dbar
rlabel m2contact -5 -98 -1 -94 3 Q
rlabel pdcontact -5 -85 -1 -81 3 D
rlabel polysilicon -10 -88 -9 -86 3 En
rlabel polysilicon -10 -145 -9 -143 3 En
rlabel metal1 -3 -176 1 -172 1 Qout
rlabel pdcontact 5 -184 9 -180 1 Vdd
rlabel ndcontact 5 -168 9 -164 5 Gnd
<< end >>
