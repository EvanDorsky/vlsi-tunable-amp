magic
tech scmos
timestamp 1259953556
<< pad >>
rect 0 0 260 260
<< end >>
