magic
tech scmos
timestamp 1259953556
<< nwell >>
rect 159 323 203 361
rect 215 323 259 361
rect 271 323 315 361
<< electrodecontact >>
rect 11 341 15 345
rect 17 341 21 345
rect 23 341 27 345
rect 29 341 33 345
rect 35 341 39 345
rect 41 341 45 345
rect 47 341 51 345
rect 11 329 15 333
rect 17 329 21 333
rect 23 329 27 333
rect 29 329 33 333
rect 35 329 39 333
rect 41 329 45 333
rect 47 329 51 333
rect 11 317 15 321
rect 17 317 21 321
rect 23 317 27 321
rect 29 317 33 321
rect 35 317 39 321
rect 41 317 45 321
rect 47 317 51 321
rect 423 341 427 345
rect 429 341 433 345
rect 435 341 439 345
rect 441 341 445 345
rect 447 341 451 345
rect 453 341 457 345
rect 459 341 463 345
rect 423 329 427 333
rect 429 329 433 333
rect 435 329 439 333
rect 441 329 445 333
rect 447 329 451 333
rect 453 329 457 333
rect 459 329 463 333
rect 423 317 427 321
rect 429 317 433 321
rect 435 317 439 321
rect 441 317 445 321
rect 447 317 451 321
rect 453 317 457 321
rect 459 317 463 321
<< electrodecap >>
rect 9 315 87 358
rect 387 315 465 358
rect 9 12 52 315
rect 422 12 465 315
<< ndiffusion >>
rect 108 359 120 360
rect 108 355 109 359
rect 113 355 115 359
rect 119 355 120 359
rect 108 353 120 355
rect 108 349 109 353
rect 113 349 115 353
rect 119 349 120 353
rect 108 347 120 349
rect 108 343 109 347
rect 113 343 115 347
rect 119 343 120 347
rect 108 341 120 343
rect 108 337 109 341
rect 113 337 115 341
rect 119 337 120 341
rect 108 335 120 337
rect 108 331 109 335
rect 113 331 115 335
rect 119 331 120 335
rect 108 329 120 331
rect 108 325 109 329
rect 113 325 115 329
rect 119 325 120 329
rect 108 324 120 325
rect 134 359 146 360
rect 134 355 135 359
rect 139 355 141 359
rect 145 355 146 359
rect 134 353 146 355
rect 134 349 135 353
rect 139 349 141 353
rect 145 349 146 353
rect 134 347 146 349
rect 134 343 135 347
rect 139 343 141 347
rect 145 343 146 347
rect 134 341 146 343
rect 134 337 135 341
rect 139 337 141 341
rect 145 337 146 341
rect 134 335 146 337
rect 134 331 135 335
rect 139 331 141 335
rect 145 331 146 335
rect 134 329 146 331
rect 134 325 135 329
rect 139 325 141 329
rect 145 325 146 329
rect 134 324 146 325
rect 328 359 340 360
rect 328 355 329 359
rect 333 355 335 359
rect 339 355 340 359
rect 328 353 340 355
rect 328 349 329 353
rect 333 349 335 353
rect 339 349 340 353
rect 328 347 340 349
rect 328 343 329 347
rect 333 343 335 347
rect 339 343 340 347
rect 328 341 340 343
rect 328 337 329 341
rect 333 337 335 341
rect 339 337 340 341
rect 328 335 340 337
rect 328 331 329 335
rect 333 331 335 335
rect 339 331 340 335
rect 328 329 340 331
rect 328 325 329 329
rect 333 325 335 329
rect 339 325 340 329
rect 328 324 340 325
rect 354 359 366 360
rect 354 355 355 359
rect 359 355 361 359
rect 365 355 366 359
rect 354 353 366 355
rect 354 349 355 353
rect 359 349 361 353
rect 365 349 366 353
rect 354 347 366 349
rect 354 343 355 347
rect 359 343 361 347
rect 365 343 366 347
rect 354 341 366 343
rect 354 337 355 341
rect 359 337 361 341
rect 365 337 366 341
rect 354 335 366 337
rect 354 331 355 335
rect 359 331 361 335
rect 365 331 366 335
rect 354 329 366 331
rect 354 325 355 329
rect 359 325 361 329
rect 365 325 366 329
rect 354 324 366 325
<< pdiffusion >>
rect 172 347 190 348
rect 172 343 173 347
rect 177 343 179 347
rect 183 343 185 347
rect 189 343 190 347
rect 172 341 190 343
rect 172 337 173 341
rect 177 337 179 341
rect 183 337 185 341
rect 189 337 190 341
rect 172 336 190 337
rect 228 347 246 348
rect 228 343 229 347
rect 233 343 235 347
rect 239 343 241 347
rect 245 343 246 347
rect 228 341 246 343
rect 228 337 229 341
rect 233 337 235 341
rect 239 337 241 341
rect 245 337 246 341
rect 228 336 246 337
rect 284 347 302 348
rect 284 343 285 347
rect 289 343 291 347
rect 295 343 297 347
rect 301 343 302 347
rect 284 341 302 343
rect 284 337 285 341
rect 289 337 291 341
rect 295 337 297 341
rect 301 337 302 341
rect 284 336 302 337
<< ndcontact >>
rect 109 355 113 359
rect 115 355 119 359
rect 109 349 113 353
rect 115 349 119 353
rect 109 343 113 347
rect 115 343 119 347
rect 109 337 113 341
rect 115 337 119 341
rect 109 331 113 335
rect 115 331 119 335
rect 109 325 113 329
rect 115 325 119 329
rect 135 355 139 359
rect 141 355 145 359
rect 135 349 139 353
rect 141 349 145 353
rect 135 343 139 347
rect 141 343 145 347
rect 135 337 139 341
rect 141 337 145 341
rect 135 331 139 335
rect 141 331 145 335
rect 135 325 139 329
rect 141 325 145 329
rect 329 355 333 359
rect 335 355 339 359
rect 329 349 333 353
rect 335 349 339 353
rect 329 343 333 347
rect 335 343 339 347
rect 329 337 333 341
rect 335 337 339 341
rect 329 331 333 335
rect 335 331 339 335
rect 329 325 333 329
rect 335 325 339 329
rect 355 355 359 359
rect 361 355 365 359
rect 355 349 359 353
rect 361 349 365 353
rect 355 343 359 347
rect 361 343 365 347
rect 355 337 359 341
rect 361 337 365 341
rect 355 331 359 335
rect 361 331 365 335
rect 355 325 359 329
rect 361 325 365 329
<< pdcontact >>
rect 173 343 177 347
rect 179 343 183 347
rect 185 343 189 347
rect 173 337 177 341
rect 179 337 183 341
rect 185 337 189 341
rect 229 343 233 347
rect 235 343 239 347
rect 241 343 245 347
rect 229 337 233 341
rect 235 337 239 341
rect 241 337 245 341
rect 285 343 289 347
rect 291 343 295 347
rect 297 343 301 347
rect 285 337 289 341
rect 291 337 295 341
rect 297 337 301 341
<< psubstratepdiff >>
rect 98 361 104 364
rect 98 357 99 361
rect 103 357 104 361
rect 124 361 130 364
rect 98 355 104 357
rect 98 351 99 355
rect 103 351 104 355
rect 98 349 104 351
rect 98 345 99 349
rect 103 345 104 349
rect 98 343 104 345
rect 98 339 99 343
rect 103 339 104 343
rect 98 337 104 339
rect 98 333 99 337
rect 103 333 104 337
rect 98 331 104 333
rect 98 327 99 331
rect 103 327 104 331
rect 98 325 104 327
rect 98 321 99 325
rect 103 321 104 325
rect 124 357 125 361
rect 129 357 130 361
rect 150 361 156 364
rect 124 355 130 357
rect 124 351 125 355
rect 129 351 130 355
rect 124 349 130 351
rect 124 345 125 349
rect 129 345 130 349
rect 124 343 130 345
rect 124 339 125 343
rect 129 339 130 343
rect 124 337 130 339
rect 124 333 125 337
rect 129 333 130 337
rect 124 331 130 333
rect 124 327 125 331
rect 129 327 130 331
rect 98 320 104 321
rect 124 320 130 327
rect 150 357 151 361
rect 155 357 156 361
rect 206 361 212 364
rect 150 355 156 357
rect 150 351 151 355
rect 155 351 156 355
rect 150 349 156 351
rect 150 345 151 349
rect 155 345 156 349
rect 150 343 156 345
rect 150 339 151 343
rect 155 339 156 343
rect 150 337 156 339
rect 150 333 151 337
rect 155 333 156 337
rect 150 331 156 333
rect 150 327 151 331
rect 155 327 156 331
rect 150 320 156 327
rect 206 357 207 361
rect 211 357 212 361
rect 262 361 268 364
rect 206 355 212 357
rect 206 351 207 355
rect 211 351 212 355
rect 206 349 212 351
rect 206 345 207 349
rect 211 345 212 349
rect 206 343 212 345
rect 206 339 207 343
rect 211 339 212 343
rect 206 337 212 339
rect 206 333 207 337
rect 211 333 212 337
rect 206 331 212 333
rect 206 327 207 331
rect 211 327 212 331
rect 206 320 212 327
rect 262 357 263 361
rect 267 357 268 361
rect 318 361 324 364
rect 262 355 268 357
rect 262 351 263 355
rect 267 351 268 355
rect 262 349 268 351
rect 262 345 263 349
rect 267 345 268 349
rect 262 343 268 345
rect 262 339 263 343
rect 267 339 268 343
rect 262 337 268 339
rect 262 333 263 337
rect 267 333 268 337
rect 262 331 268 333
rect 262 327 263 331
rect 267 327 268 331
rect 262 320 268 327
rect 318 357 319 361
rect 323 357 324 361
rect 344 361 350 364
rect 318 355 324 357
rect 318 351 319 355
rect 323 351 324 355
rect 318 349 324 351
rect 318 345 319 349
rect 323 345 324 349
rect 318 343 324 345
rect 318 339 319 343
rect 323 339 324 343
rect 318 337 324 339
rect 318 333 319 337
rect 323 333 324 337
rect 318 331 324 333
rect 318 327 319 331
rect 323 327 324 331
rect 318 320 324 327
rect 344 357 345 361
rect 349 357 350 361
rect 370 361 376 364
rect 344 355 350 357
rect 344 351 345 355
rect 349 351 350 355
rect 344 349 350 351
rect 344 345 345 349
rect 349 345 350 349
rect 344 343 350 345
rect 344 339 345 343
rect 349 339 350 343
rect 344 337 350 339
rect 344 333 345 337
rect 349 333 350 337
rect 344 331 350 333
rect 344 327 345 331
rect 349 327 350 331
rect 344 320 350 327
rect 370 357 371 361
rect 375 357 376 361
rect 370 355 376 357
rect 370 351 371 355
rect 375 351 376 355
rect 370 349 376 351
rect 370 345 371 349
rect 375 345 376 349
rect 370 343 376 345
rect 370 339 371 343
rect 375 339 376 343
rect 370 337 376 339
rect 370 333 371 337
rect 375 333 376 337
rect 370 331 376 333
rect 370 327 371 331
rect 375 327 376 331
rect 370 325 376 327
rect 370 321 371 325
rect 375 321 376 325
rect 370 320 376 321
rect 98 319 376 320
rect 98 315 99 319
rect 103 315 371 319
rect 375 315 376 319
rect 98 314 376 315
<< nsubstratendiff >>
rect 162 357 200 358
rect 162 353 163 357
rect 167 353 175 357
rect 179 353 183 357
rect 187 353 195 357
rect 199 353 200 357
rect 162 352 200 353
rect 162 349 168 352
rect 162 345 163 349
rect 167 345 168 349
rect 194 349 200 352
rect 162 341 168 345
rect 162 337 163 341
rect 167 337 168 341
rect 162 333 168 337
rect 194 345 195 349
rect 199 345 200 349
rect 194 341 200 345
rect 194 337 195 341
rect 199 337 200 341
rect 162 329 163 333
rect 167 332 168 333
rect 194 333 200 337
rect 194 332 195 333
rect 167 329 195 332
rect 199 329 200 333
rect 162 326 200 329
rect 218 357 256 358
rect 218 353 219 357
rect 223 353 251 357
rect 255 353 256 357
rect 218 352 256 353
rect 218 349 224 352
rect 218 345 219 349
rect 223 345 224 349
rect 250 349 256 352
rect 218 341 224 345
rect 218 337 219 341
rect 223 337 224 341
rect 218 333 224 337
rect 250 345 251 349
rect 255 345 256 349
rect 250 341 256 345
rect 250 337 251 341
rect 255 337 256 341
rect 218 329 219 333
rect 223 332 224 333
rect 250 333 256 337
rect 250 332 251 333
rect 223 329 251 332
rect 255 329 256 333
rect 218 326 256 329
rect 274 357 312 358
rect 274 353 275 357
rect 279 353 287 357
rect 291 353 295 357
rect 299 353 307 357
rect 311 353 312 357
rect 274 352 312 353
rect 274 349 280 352
rect 274 345 275 349
rect 279 345 280 349
rect 306 349 312 352
rect 274 341 280 345
rect 274 337 275 341
rect 279 337 280 341
rect 274 333 280 337
rect 306 345 307 349
rect 311 345 312 349
rect 306 341 312 345
rect 306 337 307 341
rect 311 337 312 341
rect 274 329 275 333
rect 279 332 280 333
rect 306 333 312 337
rect 306 332 307 333
rect 279 329 307 332
rect 311 329 312 333
rect 274 326 312 329
<< psubstratepcontact >>
rect 99 357 103 361
rect 99 351 103 355
rect 99 345 103 349
rect 99 339 103 343
rect 99 333 103 337
rect 99 327 103 331
rect 99 321 103 325
rect 125 357 129 361
rect 125 351 129 355
rect 125 345 129 349
rect 125 339 129 343
rect 125 333 129 337
rect 125 327 129 331
rect 151 357 155 361
rect 151 351 155 355
rect 151 345 155 349
rect 151 339 155 343
rect 151 333 155 337
rect 151 327 155 331
rect 207 357 211 361
rect 207 351 211 355
rect 207 345 211 349
rect 207 339 211 343
rect 207 333 211 337
rect 207 327 211 331
rect 263 357 267 361
rect 263 351 267 355
rect 263 345 267 349
rect 263 339 267 343
rect 263 333 267 337
rect 263 327 267 331
rect 319 357 323 361
rect 319 351 323 355
rect 319 345 323 349
rect 319 339 323 343
rect 319 333 323 337
rect 319 327 323 331
rect 345 357 349 361
rect 345 351 349 355
rect 345 345 349 349
rect 345 339 349 343
rect 345 333 349 337
rect 345 327 349 331
rect 371 357 375 361
rect 371 351 375 355
rect 371 345 375 349
rect 371 339 375 343
rect 371 333 375 337
rect 371 327 375 331
rect 371 321 375 325
rect 99 315 103 319
rect 371 315 375 319
<< nsubstratencontact >>
rect 163 353 167 357
rect 175 353 179 357
rect 183 353 187 357
rect 195 353 199 357
rect 163 345 167 349
rect 163 337 167 341
rect 195 345 199 349
rect 195 337 199 341
rect 163 329 167 333
rect 195 329 199 333
rect 219 353 223 357
rect 251 353 255 357
rect 219 345 223 349
rect 219 337 223 341
rect 251 345 255 349
rect 251 337 255 341
rect 219 329 223 333
rect 251 329 255 333
rect 275 353 279 357
rect 287 353 291 357
rect 295 353 299 357
rect 307 353 311 357
rect 275 345 279 349
rect 275 337 279 341
rect 307 345 311 349
rect 307 337 311 341
rect 275 329 279 333
rect 307 329 311 333
<< polysilicon >>
rect 4 361 97 363
rect 4 357 92 361
rect 96 357 97 361
rect 4 355 97 357
rect 4 351 92 355
rect 96 351 97 355
rect 4 349 97 351
rect 4 345 92 349
rect 96 345 97 349
rect 4 343 97 345
rect 4 339 92 343
rect 96 339 97 343
rect 4 337 97 339
rect 4 333 92 337
rect 96 333 97 337
rect 4 331 97 333
rect 4 327 92 331
rect 96 327 97 331
rect 4 325 97 327
rect 4 321 92 325
rect 96 321 97 325
rect 4 319 97 321
rect 4 315 92 319
rect 96 315 97 319
rect 4 310 97 315
rect 377 361 470 363
rect 377 357 378 361
rect 382 357 470 361
rect 377 355 470 357
rect 377 351 378 355
rect 382 351 470 355
rect 377 349 470 351
rect 377 345 378 349
rect 382 345 470 349
rect 377 343 470 345
rect 377 339 378 343
rect 382 339 470 343
rect 377 337 470 339
rect 377 333 378 337
rect 382 333 470 337
rect 377 331 470 333
rect 377 327 378 331
rect 382 327 470 331
rect 377 325 470 327
rect 377 321 378 325
rect 382 321 470 325
rect 377 319 470 321
rect 377 315 378 319
rect 382 315 470 319
rect 377 310 470 315
rect 4 7 57 310
rect 4 3 5 7
rect 9 3 11 7
rect 15 3 17 7
rect 21 3 23 7
rect 27 3 29 7
rect 33 3 35 7
rect 39 3 41 7
rect 45 3 47 7
rect 51 3 57 7
rect 4 2 57 3
rect 417 7 470 310
rect 417 3 423 7
rect 427 3 429 7
rect 433 3 435 7
rect 439 3 441 7
rect 445 3 447 7
rect 451 3 453 7
rect 457 3 459 7
rect 463 3 465 7
rect 469 3 470 7
rect 417 2 470 3
<< polycontact >>
rect 92 357 96 361
rect 92 351 96 355
rect 92 345 96 349
rect 92 339 96 343
rect 92 333 96 337
rect 92 327 96 331
rect 92 321 96 325
rect 92 315 96 319
rect 378 357 382 361
rect 378 351 382 355
rect 378 345 382 349
rect 378 339 382 343
rect 378 333 382 337
rect 378 327 382 331
rect 378 321 382 325
rect 378 315 382 319
rect 5 3 9 7
rect 11 3 15 7
rect 17 3 21 7
rect 23 3 27 7
rect 29 3 33 7
rect 35 3 39 7
rect 41 3 45 7
rect 47 3 51 7
rect 423 3 427 7
rect 429 3 433 7
rect 435 3 439 7
rect 441 3 445 7
rect 447 3 451 7
rect 453 3 457 7
rect 459 3 463 7
rect 465 3 469 7
<< metal1 >>
rect 229 509 230 513
rect 244 509 245 513
rect -2 365 224 369
rect -2 7 2 365
rect 99 361 103 365
rect 96 357 99 361
rect 125 361 129 365
rect 92 355 103 357
rect 96 351 99 355
rect 15 347 17 351
rect 21 347 23 351
rect 27 347 29 351
rect 33 347 35 351
rect 39 347 41 351
rect 45 347 47 351
rect 11 345 51 347
rect 15 341 17 345
rect 21 341 23 345
rect 27 341 29 345
rect 33 341 35 345
rect 39 341 41 345
rect 45 341 47 345
rect 11 339 51 341
rect 15 335 17 339
rect 21 335 23 339
rect 27 335 29 339
rect 33 335 35 339
rect 39 335 41 339
rect 45 335 47 339
rect 11 333 51 335
rect 15 329 17 333
rect 21 329 23 333
rect 27 329 29 333
rect 33 329 35 333
rect 39 329 41 333
rect 45 329 47 333
rect 11 327 51 329
rect 15 323 17 327
rect 21 323 23 327
rect 27 323 29 327
rect 33 323 35 327
rect 39 323 41 327
rect 45 323 47 327
rect 11 321 51 323
rect 15 317 17 321
rect 21 317 23 321
rect 27 317 29 321
rect 33 317 35 321
rect 39 317 41 321
rect 45 317 47 321
rect 92 349 103 351
rect 96 345 99 349
rect 92 343 103 345
rect 96 339 99 343
rect 92 337 103 339
rect 96 333 99 337
rect 92 331 103 333
rect 96 327 99 331
rect 92 325 103 327
rect 96 321 99 325
rect 92 319 103 321
rect 96 315 99 319
rect 113 355 115 359
rect 109 353 119 355
rect 113 349 115 353
rect 109 347 119 349
rect 113 343 115 347
rect 109 341 119 343
rect 113 337 115 341
rect 109 335 119 337
rect 113 331 115 335
rect 109 329 119 331
rect 113 325 115 329
rect 151 361 155 365
rect 125 355 129 357
rect 125 349 129 351
rect 125 343 129 345
rect 125 337 129 339
rect 125 331 129 333
rect 139 355 141 359
rect 135 353 145 355
rect 139 349 141 353
rect 135 347 145 349
rect 139 343 141 347
rect 135 341 145 343
rect 139 337 141 341
rect 135 335 145 337
rect 139 331 141 335
rect 135 329 145 331
rect 109 323 119 325
rect 139 325 141 329
rect 207 361 211 365
rect 151 355 155 357
rect 151 349 155 351
rect 151 343 155 345
rect 151 337 155 339
rect 151 331 155 333
rect 167 353 171 357
rect 191 353 195 357
rect 177 343 179 347
rect 183 343 185 347
rect 173 341 189 343
rect 177 337 179 341
rect 183 337 185 341
rect 135 323 145 325
rect 173 323 189 337
rect 207 355 211 357
rect 207 349 211 351
rect 207 343 211 345
rect 207 337 211 339
rect 207 331 211 333
rect 229 347 245 509
rect 250 365 476 369
rect 263 361 267 365
rect 319 361 323 365
rect 345 361 349 365
rect 233 343 235 347
rect 239 343 241 347
rect 229 341 245 343
rect 233 337 235 341
rect 239 337 241 341
rect 229 323 245 337
rect 263 355 267 357
rect 263 349 267 351
rect 263 343 267 345
rect 263 337 267 339
rect 263 331 267 333
rect 279 353 283 357
rect 303 353 307 357
rect 289 343 291 347
rect 295 343 297 347
rect 285 341 301 343
rect 289 337 291 341
rect 295 337 297 341
rect 285 323 301 337
rect 319 355 323 357
rect 319 349 323 351
rect 319 343 323 345
rect 319 337 323 339
rect 319 331 323 333
rect 333 355 335 359
rect 329 353 339 355
rect 333 349 335 353
rect 329 347 339 349
rect 333 343 335 347
rect 329 341 339 343
rect 333 337 335 341
rect 329 335 339 337
rect 333 331 335 335
rect 329 329 339 331
rect 333 325 335 329
rect 371 361 375 365
rect 345 355 349 357
rect 345 349 349 351
rect 345 343 349 345
rect 345 337 349 339
rect 345 331 349 333
rect 359 355 361 359
rect 355 353 365 355
rect 359 349 361 353
rect 355 347 365 349
rect 359 343 361 347
rect 355 341 365 343
rect 359 337 361 341
rect 355 335 365 337
rect 359 331 361 335
rect 355 329 365 331
rect 329 323 339 325
rect 359 325 361 329
rect 355 323 365 325
rect 109 310 365 323
rect 375 357 378 361
rect 371 355 382 357
rect 375 351 378 355
rect 371 349 382 351
rect 375 345 378 349
rect 371 343 382 345
rect 375 339 378 343
rect 371 337 382 339
rect 375 333 378 337
rect 371 331 382 333
rect 375 327 378 331
rect 371 325 382 327
rect 375 321 378 325
rect 371 319 382 321
rect 375 315 378 319
rect 427 347 429 351
rect 433 347 435 351
rect 439 347 441 351
rect 445 347 447 351
rect 451 347 453 351
rect 457 347 459 351
rect 423 345 463 347
rect 427 341 429 345
rect 433 341 435 345
rect 439 341 441 345
rect 445 341 447 345
rect 451 341 453 345
rect 457 341 459 345
rect 423 339 463 341
rect 427 335 429 339
rect 433 335 435 339
rect 439 335 441 339
rect 445 335 447 339
rect 451 335 453 339
rect 457 335 459 339
rect 423 333 463 335
rect 427 329 429 333
rect 433 329 435 333
rect 439 329 441 333
rect 445 329 447 333
rect 451 329 453 333
rect 457 329 459 333
rect 423 327 463 329
rect 427 323 429 327
rect 433 323 435 327
rect 439 323 441 327
rect 445 323 447 327
rect 451 323 453 327
rect 457 323 459 327
rect 423 321 463 323
rect 427 317 429 321
rect 433 317 435 321
rect 439 317 441 321
rect 445 317 447 321
rect 451 317 453 321
rect 457 317 459 321
rect 229 260 245 310
rect 472 7 476 365
rect -2 3 5 7
rect 9 3 11 7
rect 15 3 17 7
rect 21 3 23 7
rect 27 3 29 7
rect 33 3 35 7
rect 39 3 41 7
rect 45 3 47 7
rect 427 3 429 7
rect 433 3 435 7
rect 439 3 441 7
rect 445 3 447 7
rect 451 3 453 7
rect 457 3 459 7
rect 463 3 465 7
rect 469 3 476 7
<< m2contact >>
rect 230 509 244 513
rect 11 347 15 351
rect 17 347 21 351
rect 23 347 27 351
rect 29 347 33 351
rect 35 347 39 351
rect 41 347 45 351
rect 47 347 51 351
rect 11 335 15 339
rect 17 335 21 339
rect 23 335 27 339
rect 29 335 33 339
rect 35 335 39 339
rect 41 335 45 339
rect 47 335 51 339
rect 11 323 15 327
rect 17 323 21 327
rect 23 323 27 327
rect 29 323 33 327
rect 35 323 39 327
rect 41 323 45 327
rect 47 323 51 327
rect 171 353 175 357
rect 179 353 183 357
rect 187 353 191 357
rect 163 349 167 353
rect 195 349 199 353
rect 163 341 167 345
rect 163 333 167 337
rect 195 341 199 345
rect 195 333 199 337
rect 219 349 223 353
rect 219 341 223 345
rect 219 333 223 337
rect 251 349 255 353
rect 251 341 255 345
rect 251 333 255 337
rect 283 353 287 357
rect 291 353 295 357
rect 299 353 303 357
rect 275 349 279 353
rect 307 349 311 353
rect 275 341 279 345
rect 275 333 279 337
rect 307 341 311 345
rect 307 333 311 337
rect 423 347 427 351
rect 429 347 433 351
rect 435 347 439 351
rect 441 347 445 351
rect 447 347 451 351
rect 453 347 457 351
rect 459 347 463 351
rect 423 335 427 339
rect 429 335 433 339
rect 435 335 439 339
rect 441 335 445 339
rect 447 335 451 339
rect 453 335 457 339
rect 459 335 463 339
rect 423 323 427 327
rect 429 323 433 327
rect 435 323 439 327
rect 441 323 445 327
rect 447 323 451 327
rect 453 323 457 327
rect 459 323 463 327
<< metal2 >>
rect 229 509 230 513
rect 244 509 245 513
rect 11 351 51 367
rect 15 347 17 351
rect 21 347 23 351
rect 27 347 29 351
rect 33 347 35 351
rect 39 347 41 351
rect 45 347 47 351
rect 11 339 51 347
rect 15 335 17 339
rect 21 335 23 339
rect 27 335 29 339
rect 33 335 35 339
rect 39 335 41 339
rect 45 335 47 339
rect 11 327 51 335
rect 162 357 200 367
rect 162 353 171 357
rect 175 353 179 357
rect 183 353 187 357
rect 191 353 200 357
rect 162 349 163 353
rect 167 352 195 353
rect 167 349 168 352
rect 162 345 168 349
rect 162 341 163 345
rect 167 341 168 345
rect 162 337 168 341
rect 162 333 163 337
rect 167 333 168 337
rect 162 332 168 333
rect 194 349 195 352
rect 199 349 200 353
rect 194 345 200 349
rect 194 341 195 345
rect 199 341 200 345
rect 194 337 200 341
rect 194 333 195 337
rect 199 333 200 337
rect 194 332 200 333
rect 218 353 224 367
rect 218 349 219 353
rect 223 349 224 353
rect 218 345 224 349
rect 218 341 219 345
rect 223 341 224 345
rect 218 337 224 341
rect 218 333 219 337
rect 223 333 224 337
rect 218 332 224 333
rect 250 353 256 367
rect 250 349 251 353
rect 255 349 256 353
rect 250 345 256 349
rect 250 341 251 345
rect 255 341 256 345
rect 250 337 256 341
rect 250 333 251 337
rect 255 333 256 337
rect 250 332 256 333
rect 274 357 312 367
rect 274 353 283 357
rect 287 353 291 357
rect 295 353 299 357
rect 303 353 312 357
rect 274 349 275 353
rect 279 352 307 353
rect 279 349 280 352
rect 274 345 280 349
rect 274 341 275 345
rect 279 341 280 345
rect 274 337 280 341
rect 274 333 275 337
rect 279 333 280 337
rect 274 332 280 333
rect 306 349 307 352
rect 311 349 312 353
rect 306 345 312 349
rect 306 341 307 345
rect 311 341 312 345
rect 306 337 312 341
rect 306 333 307 337
rect 311 333 312 337
rect 306 332 312 333
rect 423 351 463 367
rect 427 347 429 351
rect 433 347 435 351
rect 439 347 441 351
rect 445 347 447 351
rect 451 347 453 351
rect 457 347 459 351
rect 423 339 463 347
rect 427 335 429 339
rect 433 335 435 339
rect 439 335 441 339
rect 445 335 447 339
rect 451 335 453 339
rect 457 335 459 339
rect 15 323 17 327
rect 21 323 23 327
rect 27 323 29 327
rect 33 323 35 327
rect 39 323 41 327
rect 45 323 47 327
rect 11 317 51 323
rect 423 327 463 335
rect 427 323 429 327
rect 433 323 435 327
rect 439 323 441 327
rect 445 323 447 327
rect 451 323 453 327
rect 457 323 459 327
rect 423 317 463 323
use bondingpad  bondingpad_0
timestamp 1259953556
transform 1 0 107 0 1 0
box 0 0 260 260
<< labels >>
rlabel m2contact 237 512 237 512 6 Inor
<< end >>
