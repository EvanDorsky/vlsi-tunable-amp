magic
tech scmos
timestamp 1259953556
<< electrodecontact >>
rect 11 341 15 345
rect 17 341 21 345
rect 23 341 27 345
rect 29 341 33 345
rect 35 341 39 345
rect 41 341 45 345
rect 47 341 51 345
rect 11 329 15 333
rect 17 329 21 333
rect 23 329 27 333
rect 29 329 33 333
rect 35 329 39 333
rect 41 329 45 333
rect 47 329 51 333
rect 11 317 15 321
rect 17 317 21 321
rect 23 317 27 321
rect 29 317 33 321
rect 35 317 39 321
rect 41 317 45 321
rect 47 317 51 321
rect 423 341 427 345
rect 429 341 433 345
rect 435 341 439 345
rect 441 341 445 345
rect 447 341 451 345
rect 453 341 457 345
rect 459 341 463 345
rect 423 329 427 333
rect 429 329 433 333
rect 435 329 439 333
rect 441 329 445 333
rect 447 329 451 333
rect 453 329 457 333
rect 459 329 463 333
rect 423 317 427 321
rect 429 317 433 321
rect 435 317 439 321
rect 441 317 445 321
rect 447 317 451 321
rect 453 317 457 321
rect 459 317 463 321
<< electrodecap >>
rect 9 353 123 358
rect 173 353 301 358
rect 351 353 465 358
rect 9 315 465 353
rect 9 12 52 315
rect 422 12 465 315
<< polysilicon >>
rect 4 362 470 363
rect 4 358 128 362
rect 132 358 134 362
rect 138 358 140 362
rect 144 358 146 362
rect 150 358 152 362
rect 156 358 158 362
rect 162 358 164 362
rect 168 358 306 362
rect 310 358 312 362
rect 316 358 318 362
rect 322 358 324 362
rect 328 358 330 362
rect 334 358 336 362
rect 340 358 342 362
rect 346 358 470 362
rect 4 310 470 358
rect 4 7 57 310
rect 4 3 5 7
rect 9 3 11 7
rect 15 3 17 7
rect 21 3 23 7
rect 27 3 29 7
rect 33 3 35 7
rect 39 3 41 7
rect 45 3 47 7
rect 51 3 57 7
rect 4 2 57 3
rect 417 7 470 310
rect 417 3 423 7
rect 427 3 429 7
rect 433 3 435 7
rect 439 3 441 7
rect 445 3 447 7
rect 451 3 453 7
rect 457 3 459 7
rect 463 3 465 7
rect 469 3 470 7
rect 417 2 470 3
<< polycontact >>
rect 128 358 132 362
rect 134 358 138 362
rect 140 358 144 362
rect 146 358 150 362
rect 152 358 156 362
rect 158 358 162 362
rect 164 358 168 362
rect 306 358 310 362
rect 312 358 316 362
rect 318 358 322 362
rect 324 358 328 362
rect 330 358 334 362
rect 336 358 340 362
rect 342 358 346 362
rect 5 3 9 7
rect 11 3 15 7
rect 17 3 21 7
rect 23 3 27 7
rect 29 3 33 7
rect 35 3 39 7
rect 41 3 45 7
rect 47 3 51 7
rect 423 3 427 7
rect 429 3 433 7
rect 435 3 439 7
rect 441 3 445 7
rect 447 3 451 7
rect 453 3 457 7
rect 459 3 463 7
rect 465 3 469 7
<< metal1 >>
rect 229 509 230 513
rect 244 509 245 513
rect -2 365 224 369
rect -2 7 2 365
rect 128 362 168 365
rect 132 358 134 362
rect 138 358 140 362
rect 144 358 146 362
rect 150 358 152 362
rect 156 358 158 362
rect 162 358 164 362
rect 15 347 17 351
rect 21 347 23 351
rect 27 347 29 351
rect 33 347 35 351
rect 39 347 41 351
rect 45 347 47 351
rect 11 345 51 347
rect 15 341 17 345
rect 21 341 23 345
rect 27 341 29 345
rect 33 341 35 345
rect 39 341 41 345
rect 45 341 47 345
rect 11 339 51 341
rect 15 335 17 339
rect 21 335 23 339
rect 27 335 29 339
rect 33 335 35 339
rect 39 335 41 339
rect 45 335 47 339
rect 11 333 51 335
rect 15 329 17 333
rect 21 329 23 333
rect 27 329 29 333
rect 33 329 35 333
rect 39 329 41 333
rect 45 329 47 333
rect 11 327 51 329
rect 15 323 17 327
rect 21 323 23 327
rect 27 323 29 327
rect 33 323 35 327
rect 39 323 41 327
rect 45 323 47 327
rect 11 321 51 323
rect 15 317 17 321
rect 21 317 23 321
rect 27 317 29 321
rect 33 317 35 321
rect 39 317 41 321
rect 45 317 47 321
rect 229 260 245 509
rect 250 365 476 369
rect 306 362 346 365
rect 310 358 312 362
rect 316 358 318 362
rect 322 358 324 362
rect 328 358 330 362
rect 334 358 336 362
rect 340 358 342 362
rect 427 347 429 351
rect 433 347 435 351
rect 439 347 441 351
rect 445 347 447 351
rect 451 347 453 351
rect 457 347 459 351
rect 423 345 463 347
rect 427 341 429 345
rect 433 341 435 345
rect 439 341 441 345
rect 445 341 447 345
rect 451 341 453 345
rect 457 341 459 345
rect 423 339 463 341
rect 427 335 429 339
rect 433 335 435 339
rect 439 335 441 339
rect 445 335 447 339
rect 451 335 453 339
rect 457 335 459 339
rect 423 333 463 335
rect 427 329 429 333
rect 433 329 435 333
rect 439 329 441 333
rect 445 329 447 333
rect 451 329 453 333
rect 457 329 459 333
rect 423 327 463 329
rect 427 323 429 327
rect 433 323 435 327
rect 439 323 441 327
rect 445 323 447 327
rect 451 323 453 327
rect 457 323 459 327
rect 423 321 463 323
rect 427 317 429 321
rect 433 317 435 321
rect 439 317 441 321
rect 445 317 447 321
rect 451 317 453 321
rect 457 317 459 321
rect 472 7 476 365
rect -2 3 5 7
rect 9 3 11 7
rect 15 3 17 7
rect 21 3 23 7
rect 27 3 29 7
rect 33 3 35 7
rect 39 3 41 7
rect 45 3 47 7
rect 427 3 429 7
rect 433 3 435 7
rect 439 3 441 7
rect 445 3 447 7
rect 451 3 453 7
rect 457 3 459 7
rect 463 3 465 7
rect 469 3 476 7
<< m2contact >>
rect 230 509 244 513
rect 11 347 15 351
rect 17 347 21 351
rect 23 347 27 351
rect 29 347 33 351
rect 35 347 39 351
rect 41 347 45 351
rect 47 347 51 351
rect 11 335 15 339
rect 17 335 21 339
rect 23 335 27 339
rect 29 335 33 339
rect 35 335 39 339
rect 41 335 45 339
rect 47 335 51 339
rect 11 323 15 327
rect 17 323 21 327
rect 23 323 27 327
rect 29 323 33 327
rect 35 323 39 327
rect 41 323 45 327
rect 47 323 51 327
rect 423 347 427 351
rect 429 347 433 351
rect 435 347 439 351
rect 441 347 445 351
rect 447 347 451 351
rect 453 347 457 351
rect 459 347 463 351
rect 423 335 427 339
rect 429 335 433 339
rect 435 335 439 339
rect 441 335 445 339
rect 447 335 451 339
rect 453 335 457 339
rect 459 335 463 339
rect 423 323 427 327
rect 429 323 433 327
rect 435 323 439 327
rect 441 323 445 327
rect 447 323 451 327
rect 453 323 457 327
rect 459 323 463 327
<< metal2 >>
rect 229 509 230 513
rect 244 509 245 513
rect 11 351 51 367
rect 15 347 17 351
rect 21 347 23 351
rect 27 347 29 351
rect 33 347 35 351
rect 39 347 41 351
rect 45 347 47 351
rect 11 339 51 347
rect 15 335 17 339
rect 21 335 23 339
rect 27 335 29 339
rect 33 335 35 339
rect 39 335 41 339
rect 45 335 47 339
rect 11 327 51 335
rect 15 323 17 327
rect 21 323 23 327
rect 27 323 29 327
rect 33 323 35 327
rect 39 323 41 327
rect 45 323 47 327
rect 11 317 51 323
rect 423 351 463 367
rect 427 347 429 351
rect 433 347 435 351
rect 439 347 441 351
rect 445 347 447 351
rect 451 347 453 351
rect 457 347 459 351
rect 423 339 463 347
rect 427 335 429 339
rect 433 335 435 339
rect 439 335 441 339
rect 445 335 447 339
rect 451 335 453 339
rect 457 335 459 339
rect 423 327 463 335
rect 427 323 429 327
rect 433 323 435 327
rect 439 323 441 327
rect 445 323 447 327
rect 451 323 453 327
rect 457 323 459 327
rect 423 317 463 323
use bondingpad  bondingpad_0
timestamp 1259953556
transform 1 0 107 0 1 0
box 0 0 260 260
<< labels >>
rlabel m2contact 237 512 237 512 6 Bare
<< end >>
