magic
tech scmos
timestamp 1418850683
<< nwell >>
rect 58 0 62 3
rect 43 -4 86 0
rect 142 0 146 1
rect 129 -4 172 0
rect 0 -136 2 -4
rect 58 -5 62 -4
rect 153 -5 157 -4
<< pwell >>
rect 0 -4 43 3
rect 86 -4 129 3
rect 0 -388 2 -136
<< electrodecontact >>
rect 1084 -9 1088 141
<< electrodecap >>
rect 1082 -13 1238 143
<< ptransistor >>
rect 296 -11 302 229
rect 308 -11 314 229
rect 320 -11 326 229
rect 332 -11 338 229
rect 344 -11 350 229
rect 356 -11 362 229
rect 368 -11 374 229
rect 380 -11 386 229
rect 392 -11 398 229
rect 404 -11 410 229
rect 416 -11 422 229
rect 428 -11 434 229
rect 440 -11 446 229
rect 452 -11 458 229
rect 464 -11 470 229
rect 476 -11 482 229
rect 488 -11 494 229
rect 500 -11 506 229
rect 512 -11 518 229
rect 524 -11 530 229
rect 536 -11 542 229
rect 548 -11 554 229
rect 560 -11 566 229
rect 572 -11 578 229
rect 584 -11 590 229
rect 596 -11 602 229
rect 608 -11 614 229
rect 620 -11 626 229
rect 632 -11 638 229
rect 644 -11 650 229
rect 656 -11 662 229
rect 668 -11 674 229
rect 680 -11 686 229
rect 692 -11 698 229
rect 704 -11 710 229
rect 716 -11 722 229
rect 728 -11 734 229
rect 740 -11 746 229
rect 752 -11 758 229
rect 764 -11 770 229
rect 776 -11 782 229
rect 788 -11 794 229
rect 800 -11 806 229
rect 812 -11 818 229
rect 824 -11 830 229
rect 836 -11 842 229
rect 848 -11 854 229
rect 860 -11 866 229
rect 872 -11 878 229
rect 884 -11 890 229
<< pdiffusion >>
rect 290 -11 291 229
rect 295 -11 296 229
rect 302 -11 303 229
rect 307 -11 308 229
rect 314 -11 315 229
rect 319 -11 320 229
rect 326 -11 327 229
rect 331 -11 332 229
rect 338 -11 339 229
rect 343 -11 344 229
rect 350 -11 351 229
rect 355 -11 356 229
rect 362 -11 363 229
rect 367 -11 368 229
rect 374 -11 375 229
rect 379 -11 380 229
rect 386 -11 387 229
rect 391 -11 392 229
rect 398 -11 399 229
rect 403 -11 404 229
rect 410 -11 411 229
rect 415 -11 416 229
rect 422 -11 423 229
rect 427 -11 428 229
rect 434 -11 435 229
rect 439 -11 440 229
rect 446 -11 447 229
rect 451 -11 452 229
rect 458 -11 459 229
rect 463 -11 464 229
rect 470 -11 471 229
rect 475 -11 476 229
rect 482 -11 483 229
rect 487 -11 488 229
rect 494 -11 495 229
rect 499 -11 500 229
rect 506 -11 507 229
rect 511 -11 512 229
rect 518 -11 519 229
rect 523 -11 524 229
rect 530 -11 531 229
rect 535 -11 536 229
rect 542 -11 543 229
rect 547 -11 548 229
rect 554 -11 555 229
rect 559 -11 560 229
rect 566 -11 567 229
rect 571 -11 572 229
rect 578 -11 579 229
rect 583 -11 584 229
rect 590 -11 591 229
rect 595 -11 596 229
rect 602 -11 603 229
rect 607 -11 608 229
rect 614 -11 615 229
rect 619 -11 620 229
rect 626 -11 627 229
rect 631 -11 632 229
rect 638 -11 639 229
rect 643 -11 644 229
rect 650 -11 651 229
rect 655 -11 656 229
rect 662 -11 663 229
rect 667 -11 668 229
rect 674 -11 675 229
rect 679 -11 680 229
rect 686 -11 687 229
rect 691 -11 692 229
rect 698 -11 699 229
rect 703 -11 704 229
rect 710 -11 711 229
rect 715 -11 716 229
rect 722 -11 723 229
rect 727 -11 728 229
rect 734 -11 735 229
rect 739 -11 740 229
rect 746 -11 747 229
rect 751 -11 752 229
rect 758 -11 759 229
rect 763 -11 764 229
rect 770 -11 771 229
rect 775 -11 776 229
rect 782 -11 783 229
rect 787 -11 788 229
rect 794 -11 795 229
rect 799 -11 800 229
rect 806 -11 807 229
rect 811 -11 812 229
rect 818 -11 819 229
rect 823 -11 824 229
rect 830 -11 831 229
rect 835 -11 836 229
rect 842 -11 843 229
rect 847 -11 848 229
rect 854 -11 855 229
rect 859 -11 860 229
rect 866 -11 867 229
rect 871 -11 872 229
rect 878 -11 879 229
rect 883 -11 884 229
rect 890 -11 891 229
rect 895 -11 896 229
<< pdcontact >>
rect 11 -14 15 -10
rect 103 -14 107 -10
rect 291 -11 295 229
rect 303 -11 307 229
rect 315 -11 319 229
rect 327 -11 331 229
rect 339 -11 343 229
rect 351 -11 355 229
rect 363 -11 367 229
rect 375 -11 379 229
rect 387 -11 391 229
rect 399 -11 403 229
rect 411 -11 415 229
rect 423 -11 427 229
rect 435 -11 439 229
rect 447 -11 451 229
rect 459 -11 463 229
rect 471 -11 475 229
rect 483 -11 487 229
rect 495 -11 499 229
rect 507 -11 511 229
rect 519 -11 523 229
rect 531 -11 535 229
rect 543 -11 547 229
rect 555 -11 559 229
rect 567 -11 571 229
rect 579 -11 583 229
rect 591 -11 595 229
rect 603 -11 607 229
rect 615 -11 619 229
rect 627 -11 631 229
rect 639 -11 643 229
rect 651 -11 655 229
rect 663 -11 667 229
rect 675 -11 679 229
rect 687 -11 691 229
rect 699 -11 703 229
rect 711 -11 715 229
rect 723 -11 727 229
rect 735 -11 739 229
rect 747 -11 751 229
rect 759 -11 763 229
rect 771 -11 775 229
rect 783 -11 787 229
rect 795 -11 799 229
rect 807 -11 811 229
rect 819 -11 823 229
rect 831 -11 835 229
rect 843 -11 847 229
rect 855 -11 859 229
rect 867 -11 871 229
rect 879 -11 883 229
rect 891 -11 895 229
<< polysilicon >>
rect 296 229 302 232
rect 308 229 314 232
rect 320 229 326 232
rect 332 229 338 232
rect 344 229 350 232
rect 356 229 362 232
rect 368 229 374 232
rect 380 229 386 232
rect 392 229 398 232
rect 404 229 410 232
rect 416 229 422 232
rect 428 229 434 232
rect 440 229 446 232
rect 452 229 458 232
rect 464 229 470 232
rect 476 229 482 232
rect 488 229 494 232
rect 500 229 506 232
rect 512 229 518 232
rect 524 229 530 232
rect 536 229 542 232
rect 548 229 554 232
rect 560 229 566 232
rect 572 229 578 232
rect 584 229 590 232
rect 596 229 602 232
rect 608 229 614 232
rect 620 229 626 232
rect 632 229 638 232
rect 644 229 650 232
rect 656 229 662 232
rect 668 229 674 232
rect 680 229 686 232
rect 692 229 698 232
rect 704 229 710 232
rect 716 229 722 232
rect 728 229 734 232
rect 740 229 746 232
rect 752 229 758 232
rect 764 229 770 232
rect 776 229 782 232
rect 788 229 794 232
rect 800 229 806 232
rect 812 229 818 232
rect 824 229 830 232
rect 836 229 842 232
rect 848 229 854 232
rect 860 229 866 232
rect 872 229 878 232
rect 884 229 890 232
rect 57 3 63 4
rect 109 3 115 4
rect 296 -14 302 -11
rect 308 -14 314 -11
rect 320 -14 326 -11
rect 332 -14 338 -11
rect 344 -14 350 -11
rect 356 -14 362 -11
rect 368 -14 374 -11
rect 380 -14 386 -11
rect 392 -14 398 -11
rect 404 -14 410 -11
rect 416 -14 422 -11
rect 428 -14 434 -11
rect 440 -14 446 -11
rect 452 -14 458 -11
rect 464 -14 470 -11
rect 476 -14 482 -11
rect 488 -14 494 -11
rect 500 -14 506 -11
rect 512 -14 518 -11
rect 524 -14 530 -11
rect 536 -14 542 -11
rect 548 -14 554 -11
rect 560 -14 566 -11
rect 572 -14 578 -11
rect 584 -14 590 -11
rect 596 -14 602 -11
rect 608 -14 614 -11
rect 620 -14 626 -11
rect 632 -14 638 -11
rect 644 -14 650 -11
rect 656 -14 662 -11
rect 668 -14 674 -11
rect 680 -14 686 -11
rect 692 -14 698 -11
rect 704 -14 710 -11
rect 716 -14 722 -11
rect 728 -14 734 -11
rect 740 -14 746 -11
rect 752 -14 758 -11
rect 764 -14 770 -11
rect 776 -14 782 -11
rect 788 -14 794 -11
rect 800 -14 806 -11
rect 812 -14 818 -11
rect 824 -14 830 -11
rect 836 -14 842 -11
rect 848 -14 854 -11
rect 860 -14 866 -11
rect 872 -14 878 -11
rect 884 -14 890 -11
rect 290 -18 890 -14
rect 1077 -18 1243 148
<< polycontact >>
rect 26 1 30 5
rect 58 -1 62 3
rect 110 -1 114 3
rect 142 1 146 5
rect 153 -9 157 -5
<< metal1 >>
rect 293 232 890 236
rect 303 229 307 232
rect 327 229 331 232
rect 351 229 355 232
rect 375 229 379 232
rect 399 229 403 232
rect 423 229 427 232
rect 447 229 451 232
rect 471 229 475 232
rect 495 229 499 232
rect 519 229 523 232
rect 543 229 547 232
rect 567 229 571 232
rect 591 229 595 232
rect 615 229 619 232
rect 639 229 643 232
rect 663 229 667 232
rect 687 229 691 232
rect 711 229 715 232
rect 735 229 739 232
rect 759 229 763 232
rect 783 229 787 232
rect 807 229 811 232
rect 831 229 835 232
rect 855 229 859 232
rect 879 229 883 232
rect 26 -1 30 1
rect 11 -5 30 -1
rect 58 -5 62 -1
rect 103 -5 114 -1
rect 142 0 146 1
rect 142 -4 157 0
rect 153 -5 157 -4
rect 11 -10 15 -5
rect 103 -10 107 -5
rect 291 -14 295 -11
rect 315 -14 319 -11
rect 339 -14 343 -11
rect 363 -14 367 -11
rect 387 -14 391 -11
rect 411 -14 415 -11
rect 435 -14 439 -11
rect 459 -14 463 -11
rect 483 -14 487 -11
rect 507 -14 511 -11
rect 531 -14 535 -11
rect 555 -14 559 -11
rect 579 -14 583 -11
rect 603 -14 607 -11
rect 627 -14 631 -11
rect 651 -14 655 -11
rect 675 -14 679 -11
rect 699 -14 703 -11
rect 723 -14 727 -11
rect 747 -14 751 -11
rect 771 -14 775 -11
rect 795 -14 799 -11
rect 819 -14 823 -11
rect 843 -14 847 -11
rect 867 -14 871 -11
rect 891 -14 895 -11
rect 1084 -14 1088 -9
rect 290 -18 895 -14
rect 1077 -18 1088 -14
use amp  amp_0
timestamp 1418768421
transform 1 0 95 0 1 135
box -95 -135 77 126
use bias  bias_0
timestamp 1418768461
transform 1 0 -11 0 1 -106
box 13 -282 183 102
<< end >>
