magic
tech scmos
timestamp 1419261862
<< nwell >>
rect 766 603 770 607
rect 766 599 769 600
rect 766 579 770 583
rect 518 511 562 514
rect 636 511 670 514
<< pwell >>
rect 259 668 1252 698
rect 553 648 585 668
rect 753 618 756 619
rect 761 613 762 614
rect 759 612 762 613
rect 759 611 761 612
rect 760 608 761 611
rect 752 604 753 607
rect 760 597 763 608
<< electrodecontact >>
rect 1686 268 1690 420
<< psubstratepcontact >>
rect 500 671 860 675
<< polycontact >>
rect 865 518 869 522
<< metal1 >>
rect 883 691 885 692
rect 865 688 885 691
rect 266 654 269 669
rect 567 662 571 671
rect 865 668 869 688
rect 838 661 862 664
rect 1238 661 1242 669
rect 762 659 1242 661
rect 762 657 844 659
rect 858 657 1242 659
rect 545 654 593 655
rect 266 652 775 654
rect 266 651 548 652
rect 590 651 771 652
rect 753 618 756 619
rect 735 520 790 524
rect 1686 420 1689 674
<< m2contact >>
rect 480 664 484 668
rect 889 673 893 677
rect 865 664 869 668
rect 1238 669 1242 673
rect 567 658 571 662
rect 758 657 762 661
rect 567 645 571 649
rect 771 648 775 652
rect 823 625 827 629
rect 766 603 770 607
rect 766 579 770 583
rect 766 555 770 559
rect 766 531 770 535
rect 865 522 869 526
<< metal2 >>
rect 765 673 889 674
rect 765 671 892 673
rect 561 667 577 668
rect 484 665 749 667
rect 484 664 564 665
rect 574 664 749 665
rect 567 649 571 658
rect 746 636 749 664
rect 746 633 756 636
rect 753 607 756 633
rect 759 614 762 657
rect 765 620 768 671
rect 771 626 774 648
rect 777 629 786 633
rect 771 623 776 626
rect 782 625 823 629
rect 765 617 770 620
rect 759 611 763 614
rect 752 604 756 607
rect 752 576 755 604
rect 760 600 763 611
rect 767 607 770 617
rect 760 597 769 600
rect 766 583 769 597
rect 752 573 769 576
rect 766 559 769 573
rect 773 535 776 623
rect 770 532 776 535
rect 865 526 869 664
use resistors  resistors_0
timestamp 1419231588
transform -1 0 1688 0 -1 699
box -11 -21 1656 35
use spi-interface  spi-interface_0
timestamp 1418856619
transform 0 1 502 -1 0 622
box -27 -21 108 279
use amplifier  amplifier_0
timestamp 1418878488
transform 1 0 781 0 1 394
box -781 -394 952 261
<< labels >>
rlabel metal2 765 634 768 636 1 B0
rlabel metal2 759 634 762 636 1 B1
rlabel metal2 753 634 756 636 1 B2
rlabel metal2 771 634 774 636 1 B3
<< end >>
