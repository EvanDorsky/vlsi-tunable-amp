magic
tech scmos
magscale 1 3
timestamp 1419065237
<< metal1 >>
rect 2626 7276 2676 7286
rect 2596 7266 2706 7276
rect 2586 7256 2716 7266
rect 2556 7236 2716 7256
rect 2876 7236 2946 7256
rect 2536 7226 2716 7236
rect 2866 7226 2946 7236
rect 2516 7216 2706 7226
rect 2866 7216 2956 7226
rect 2976 7216 2996 7226
rect 3016 7216 3096 7226
rect 2506 7206 2686 7216
rect 2856 7206 3146 7216
rect 2486 7196 2686 7206
rect 2846 7196 3176 7206
rect 2476 7186 2666 7196
rect 2846 7186 3196 7196
rect 2446 7176 2676 7186
rect 2746 7176 2776 7186
rect 2786 7176 2806 7186
rect 2846 7176 3236 7186
rect 2436 7166 2686 7176
rect 2746 7166 2826 7176
rect 2886 7166 3246 7176
rect 2416 7156 2696 7166
rect 2726 7156 2856 7166
rect 2896 7156 3276 7166
rect 2376 7146 2866 7156
rect 2896 7146 3296 7156
rect 2366 7136 2876 7146
rect 2886 7136 2946 7146
rect 3016 7136 3036 7146
rect 3166 7136 3276 7146
rect 2346 7126 2936 7136
rect 3196 7126 3216 7136
rect 2316 7116 2926 7126
rect 2286 7106 2936 7116
rect 2266 7096 2956 7106
rect 2246 7086 2966 7096
rect 2236 7076 2966 7086
rect 2226 7066 2906 7076
rect 2926 7066 2956 7076
rect 2206 7056 2906 7066
rect 2196 7046 2906 7056
rect 2186 7036 2926 7046
rect 2176 7026 2916 7036
rect 2166 7006 2916 7026
rect 2156 6996 2916 7006
rect 2156 6986 2906 6996
rect 2146 6976 2896 6986
rect 3116 6976 3126 6996
rect 2136 6966 2736 6976
rect 2826 6966 2906 6976
rect 2116 6956 2746 6966
rect 2846 6956 2856 6966
rect 2876 6956 2896 6966
rect 2106 6946 2756 6956
rect 2106 6936 2686 6946
rect 2706 6936 2716 6946
rect 2726 6936 2756 6946
rect 3116 6946 3176 6956
rect 3116 6936 3206 6946
rect 2086 6926 2646 6936
rect 3126 6926 3266 6936
rect 2086 6916 2636 6926
rect 3156 6916 3276 6926
rect 2066 6906 2646 6916
rect 3196 6906 3306 6916
rect 2046 6896 2666 6906
rect 3236 6896 3316 6906
rect 2026 6886 2686 6896
rect 3256 6886 3326 6896
rect 2006 6876 2686 6886
rect 3286 6876 3306 6886
rect 1996 6866 2716 6876
rect 1976 6856 2736 6866
rect 1966 6846 2496 6856
rect 2586 6846 2746 6856
rect 1946 6836 2496 6846
rect 2596 6836 2756 6846
rect 1946 6826 2536 6836
rect 2606 6826 2796 6836
rect 1936 6816 2556 6826
rect 2566 6816 2586 6826
rect 2606 6816 2806 6826
rect 1946 6806 2826 6816
rect 1946 6796 2846 6806
rect 1946 6786 2896 6796
rect 1946 6776 2906 6786
rect 1946 6766 2916 6776
rect 1926 6756 2926 6766
rect 1916 6746 2596 6756
rect 2626 6746 2926 6756
rect 1906 6736 2566 6746
rect 2636 6736 2876 6746
rect 1896 6716 2566 6736
rect 2706 6726 2876 6736
rect 2726 6716 2856 6726
rect 1886 6706 2576 6716
rect 2746 6706 2856 6716
rect 1876 6696 2586 6706
rect 2786 6696 2856 6706
rect 1866 6686 2586 6696
rect 2806 6686 2866 6696
rect 3666 6686 3686 6696
rect 1846 6666 2516 6686
rect 2526 6676 2586 6686
rect 2836 6676 2886 6686
rect 3666 6676 3716 6686
rect 2536 6666 2586 6676
rect 2846 6666 2886 6676
rect 3676 6666 3716 6676
rect 1846 6656 2506 6666
rect 2566 6656 2586 6666
rect 2866 6656 2886 6666
rect 3666 6656 3766 6666
rect 1826 6636 2496 6656
rect 3626 6646 3766 6656
rect 3626 6636 3806 6646
rect 1846 6626 2176 6636
rect 2216 6626 2506 6636
rect 3646 6626 3826 6636
rect 1846 6616 2166 6626
rect 1816 6606 2156 6616
rect 2226 6606 2506 6626
rect 2966 6616 3016 6626
rect 3656 6616 3836 6626
rect 2966 6606 3026 6616
rect 3676 6606 3836 6616
rect 1816 6596 2086 6606
rect 2096 6596 2156 6606
rect 1816 6576 2156 6596
rect 1806 6566 2156 6576
rect 2196 6566 2206 6576
rect 1726 6556 1736 6566
rect 1796 6556 2156 6566
rect 2186 6556 2206 6566
rect 2236 6566 2506 6606
rect 2976 6596 3036 6606
rect 3236 6596 3276 6606
rect 3676 6596 3866 6606
rect 3006 6586 3046 6596
rect 3016 6576 3056 6586
rect 3236 6576 3296 6596
rect 3356 6586 3366 6596
rect 3396 6586 3416 6596
rect 3686 6586 3876 6596
rect 3386 6576 3436 6586
rect 3706 6576 3886 6586
rect 3036 6566 3046 6576
rect 2236 6556 2516 6566
rect 3246 6556 3286 6576
rect 3376 6566 3446 6576
rect 3706 6566 3926 6576
rect 3376 6556 3466 6566
rect 3736 6556 3926 6566
rect 1716 6546 1746 6556
rect 1796 6546 2154 6556
rect 2196 6546 2206 6556
rect 1706 6536 1756 6546
rect 1796 6536 2136 6546
rect 2246 6536 2526 6556
rect 3246 6546 3296 6556
rect 3376 6546 3406 6556
rect 3416 6546 3486 6556
rect 3746 6546 3936 6556
rect 3256 6536 3306 6546
rect 3426 6536 3506 6546
rect 3766 6536 3966 6546
rect 1706 6526 1766 6536
rect 1786 6526 2146 6536
rect 2246 6526 2536 6536
rect 3276 6526 3316 6536
rect 3436 6526 3516 6536
rect 3776 6526 3986 6536
rect 1706 6516 2146 6526
rect 2236 6516 2356 6526
rect 2386 6516 2556 6526
rect 3286 6516 3326 6526
rect 3456 6516 3536 6526
rect 3786 6516 3996 6526
rect 1696 6506 2146 6516
rect 2246 6506 2346 6516
rect 2386 6506 2566 6516
rect 1696 6496 2026 6506
rect 1686 6486 1986 6496
rect 2006 6486 2026 6496
rect 1676 6476 1936 6486
rect 1956 6476 1986 6486
rect 1666 6466 1936 6476
rect 1966 6466 1986 6476
rect 2016 6466 2026 6486
rect 2046 6476 2136 6506
rect 2246 6496 2336 6506
rect 2376 6496 2566 6506
rect 3306 6506 3326 6516
rect 3466 6506 3546 6516
rect 3796 6506 4016 6516
rect 3306 6496 3336 6506
rect 3476 6496 3546 6506
rect 3806 6496 4036 6506
rect 2256 6486 2326 6496
rect 2366 6486 2546 6496
rect 3326 6486 3366 6496
rect 3476 6486 3526 6496
rect 3816 6486 4066 6496
rect 2226 6476 2236 6486
rect 2256 6476 2316 6486
rect 2356 6476 2426 6486
rect 2056 6466 2136 6476
rect 2216 6466 2236 6476
rect 2246 6466 2306 6476
rect 2346 6466 2416 6476
rect 1656 6456 1936 6466
rect 2056 6456 2126 6466
rect 2246 6456 2296 6466
rect 1646 6436 1936 6456
rect 1636 6426 1666 6436
rect 1676 6426 1936 6436
rect 2066 6426 2126 6456
rect 2236 6446 2296 6456
rect 2336 6456 2396 6466
rect 2436 6456 2516 6486
rect 3336 6476 3376 6486
rect 3486 6476 3516 6486
rect 3826 6476 4086 6486
rect 3346 6466 3386 6476
rect 3506 6466 3556 6476
rect 3826 6466 4106 6476
rect 3356 6456 3396 6466
rect 2336 6446 2376 6456
rect 2426 6446 2526 6456
rect 3366 6446 3406 6456
rect 3516 6446 3566 6466
rect 3826 6456 4126 6466
rect 3576 6446 3586 6456
rect 3866 6446 4126 6456
rect 2236 6436 2286 6446
rect 2306 6436 2316 6446
rect 2346 6436 2356 6446
rect 2226 6426 2276 6436
rect 1636 6416 1656 6426
rect 1686 6416 1926 6426
rect 1616 6396 1626 6406
rect 1696 6396 1916 6416
rect 2066 6406 2116 6426
rect 2216 6416 2266 6426
rect 1606 6376 1626 6396
rect 1706 6386 1906 6396
rect 1716 6376 1906 6386
rect 2066 6376 2106 6406
rect 2216 6396 2276 6416
rect 2306 6406 2326 6436
rect 2416 6426 2526 6446
rect 3376 6436 3426 6446
rect 3526 6436 3536 6446
rect 3376 6426 3446 6436
rect 3546 6426 3596 6446
rect 3856 6436 4156 6446
rect 3876 6426 4166 6436
rect 2416 6416 2536 6426
rect 2406 6406 2546 6416
rect 2656 6406 2686 6426
rect 3386 6416 3456 6426
rect 3546 6416 3616 6426
rect 3886 6416 4176 6426
rect 3386 6406 3476 6416
rect 3576 6406 3616 6416
rect 3896 6406 4176 6416
rect 2406 6396 2556 6406
rect 2656 6396 2696 6406
rect 3396 6396 3476 6406
rect 3586 6396 3616 6406
rect 3906 6396 4186 6406
rect 2226 6386 2276 6396
rect 2416 6386 2566 6396
rect 2226 6376 2266 6386
rect 2406 6376 2566 6386
rect 2676 6386 2706 6396
rect 3236 6386 3256 6396
rect 3406 6386 3486 6396
rect 3676 6386 3706 6396
rect 3916 6386 4196 6396
rect 2676 6376 2726 6386
rect 3236 6376 3276 6386
rect 3426 6376 3496 6386
rect 3676 6376 3726 6386
rect 3926 6376 4196 6386
rect 1596 6366 1626 6376
rect 1726 6366 1896 6376
rect 2076 6366 2096 6376
rect 2196 6366 2256 6376
rect 2396 6366 2566 6376
rect 2686 6366 2736 6376
rect 3116 6366 3156 6376
rect 3236 6366 3296 6376
rect 1596 6356 1616 6366
rect 1726 6356 1766 6366
rect 1776 6356 1886 6366
rect 2176 6356 2236 6366
rect 2386 6356 2577 6366
rect 2726 6356 2796 6366
rect 2816 6356 2846 6366
rect 2916 6356 2936 6366
rect 3116 6356 3166 6366
rect 3216 6356 3296 6366
rect 3436 6366 3546 6376
rect 3676 6366 3776 6376
rect 3936 6366 4206 6376
rect 3436 6356 3556 6366
rect 3676 6356 3786 6366
rect 3966 6356 4206 6366
rect 1656 6346 1676 6356
rect 1726 6346 1756 6356
rect 1776 6346 1876 6356
rect 2176 6346 2226 6356
rect 2376 6346 2606 6356
rect 2736 6346 2856 6356
rect 2916 6346 2966 6356
rect 3126 6346 3316 6356
rect 3446 6346 3566 6356
rect 3686 6346 3796 6356
rect 3976 6346 4236 6356
rect 1656 6326 1686 6346
rect 1666 6316 1686 6326
rect 1776 6336 1866 6346
rect 2176 6336 2196 6346
rect 2216 6336 2226 6346
rect 2366 6336 2606 6346
rect 2746 6336 2866 6346
rect 2926 6336 2976 6346
rect 3126 6336 3156 6346
rect 3166 6336 3326 6346
rect 3456 6336 3586 6346
rect 3696 6336 3806 6346
rect 3976 6336 4286 6346
rect 1776 6316 1856 6336
rect 2366 6326 2616 6336
rect 2756 6326 2876 6336
rect 2926 6326 2986 6336
rect 3126 6326 3346 6336
rect 3466 6326 3596 6336
rect 3706 6326 3816 6336
rect 3986 6326 4296 6336
rect 2166 6316 2176 6326
rect 2366 6316 2476 6326
rect 1766 6296 1856 6316
rect 1586 6276 1606 6286
rect 1676 6276 1686 6286
rect 1586 6246 1616 6276
rect 1666 6266 1686 6276
rect 1756 6276 1846 6296
rect 2146 6286 2176 6316
rect 2256 6296 2266 6316
rect 2356 6306 2466 6316
rect 2346 6286 2466 6306
rect 2486 6296 2626 6326
rect 2766 6316 2876 6326
rect 2936 6316 3006 6326
rect 3126 6316 3366 6326
rect 3486 6316 3616 6326
rect 3716 6316 3836 6326
rect 2786 6306 2886 6316
rect 2946 6306 3006 6316
rect 3146 6306 3156 6316
rect 3166 6306 3376 6316
rect 3496 6306 3626 6316
rect 3736 6306 3846 6316
rect 3996 6306 4256 6326
rect 4276 6316 4316 6326
rect 4286 6306 4326 6316
rect 2796 6296 2896 6306
rect 2956 6296 3036 6306
rect 3146 6296 3396 6306
rect 3506 6296 3636 6306
rect 3746 6296 3856 6306
rect 4006 6296 4316 6306
rect 2146 6276 2166 6286
rect 2336 6276 2466 6286
rect 1756 6256 1836 6276
rect 2336 6266 2456 6276
rect 2326 6256 2346 6266
rect 1756 6246 1826 6256
rect 2316 6246 2346 6256
rect 1596 6226 1626 6246
rect 1756 6236 1816 6246
rect 1666 6226 1676 6236
rect 1746 6226 1806 6236
rect 2116 6226 2126 6246
rect 2316 6226 2336 6246
rect 2366 6226 2456 6266
rect 2476 6266 2656 6296
rect 2816 6286 2906 6296
rect 2966 6286 3056 6296
rect 2826 6276 2906 6286
rect 2976 6276 3056 6286
rect 3136 6286 3406 6296
rect 3506 6286 3646 6296
rect 3746 6286 3866 6296
rect 4026 6286 4326 6296
rect 3136 6276 3416 6286
rect 3506 6276 3666 6286
rect 3756 6276 3876 6286
rect 3966 6276 3976 6286
rect 4046 6276 4326 6286
rect 2836 6266 2916 6276
rect 2986 6266 3076 6276
rect 3096 6266 3106 6276
rect 3126 6266 3426 6276
rect 3516 6266 3686 6276
rect 3766 6266 3926 6276
rect 3936 6266 3986 6276
rect 4086 6266 4336 6276
rect 2476 6256 2666 6266
rect 2846 6256 2916 6266
rect 3016 6256 3446 6266
rect 3526 6256 3686 6266
rect 3776 6256 3986 6266
rect 4096 6256 4346 6266
rect 2476 6246 2676 6256
rect 2856 6246 2906 6256
rect 3026 6246 3466 6256
rect 3536 6246 3706 6256
rect 3786 6246 3996 6256
rect 4086 6246 4346 6256
rect 2476 6226 2636 6246
rect 2656 6236 2676 6246
rect 3046 6236 3466 6246
rect 3546 6236 3716 6246
rect 3796 6236 4006 6246
rect 4076 6236 4336 6246
rect 1586 6216 1676 6226
rect 1576 6206 1666 6216
rect 1736 6206 1796 6226
rect 2316 6216 2326 6226
rect 2356 6206 2446 6226
rect 1576 6196 1656 6206
rect 1586 6186 1656 6196
rect 1736 6186 1786 6206
rect 2146 6196 2156 6206
rect 2346 6196 2446 6206
rect 2126 6186 2136 6196
rect 2146 6186 2166 6196
rect 1576 6176 1666 6186
rect 1716 6176 1776 6186
rect 2116 6176 2136 6186
rect 1576 6156 1676 6176
rect 1706 6166 1766 6176
rect 1696 6156 1736 6166
rect 2286 6156 2306 6186
rect 1576 6146 1726 6156
rect 2276 6146 2306 6156
rect 2336 6176 2376 6196
rect 2406 6186 2446 6196
rect 2476 6216 2646 6226
rect 2656 6216 2686 6236
rect 3046 6226 3186 6236
rect 3216 6226 3476 6236
rect 3556 6226 3716 6236
rect 3806 6226 4026 6236
rect 4086 6226 4106 6236
rect 4126 6226 4336 6236
rect 3056 6216 3196 6226
rect 3226 6216 3476 6226
rect 3576 6216 3736 6226
rect 3816 6216 3846 6226
rect 3906 6216 4026 6226
rect 2476 6206 2696 6216
rect 3046 6206 3076 6216
rect 3086 6206 3206 6216
rect 3236 6206 3476 6216
rect 3586 6206 3746 6216
rect 3856 6206 3876 6216
rect 3896 6206 4056 6216
rect 4176 6206 4336 6226
rect 2476 6196 2706 6206
rect 3046 6196 3066 6206
rect 3106 6196 3216 6206
rect 3246 6196 3486 6206
rect 3606 6196 3756 6206
rect 3836 6196 4076 6206
rect 4186 6196 4346 6206
rect 2476 6186 2526 6196
rect 2556 6186 2716 6196
rect 3048 6195 3226 6196
rect 2406 6176 2436 6186
rect 2476 6176 2516 6186
rect 2336 6156 2366 6176
rect 2406 6166 2426 6176
rect 2396 6156 2426 6166
rect 2476 6156 2496 6176
rect 2546 6166 2716 6186
rect 3056 6186 3226 6195
rect 3256 6186 3486 6196
rect 3626 6186 3766 6196
rect 3836 6186 4096 6196
rect 4196 6186 4376 6196
rect 3056 6176 3236 6186
rect 3266 6176 3506 6186
rect 3636 6176 3806 6186
rect 3836 6176 4106 6186
rect 4216 6176 4376 6186
rect 2536 6165 2716 6166
rect 2526 6156 2716 6165
rect 3046 6166 3246 6176
rect 3286 6166 3536 6176
rect 3636 6166 3816 6176
rect 3846 6166 4106 6176
rect 4246 6166 4376 6176
rect 3046 6156 3256 6166
rect 3306 6156 3546 6166
rect 3646 6156 3826 6166
rect 3856 6156 4126 6166
rect 4246 6156 4386 6166
rect 2336 6146 2356 6156
rect 2386 6146 2416 6156
rect 2506 6153 2726 6156
rect 2506 6146 2536 6153
rect 2556 6146 2726 6153
rect 3056 6146 3296 6156
rect 1566 6136 1686 6146
rect 1556 6126 1686 6136
rect 1546 6116 1676 6126
rect 1536 6106 1676 6116
rect 1536 6066 1716 6106
rect 2266 6096 2296 6146
rect 2326 6136 2346 6146
rect 2386 6136 2406 6146
rect 2506 6136 2526 6146
rect 2556 6136 2736 6146
rect 3066 6136 3296 6146
rect 3316 6136 3546 6156
rect 3666 6146 3846 6156
rect 3856 6147 4146 6156
rect 3856 6146 4158 6147
rect 3676 6136 4158 6146
rect 4246 6146 4396 6156
rect 4246 6136 4296 6146
rect 4336 6136 4406 6146
rect 2316 6116 2346 6136
rect 2496 6116 2516 6136
rect 2266 6076 2286 6096
rect 2316 6086 2336 6116
rect 2506 6106 2516 6116
rect 2566 6126 2746 6136
rect 3076 6126 3306 6136
rect 3316 6126 3576 6136
rect 3686 6126 4126 6136
rect 4137 6135 4166 6136
rect 4146 6126 4166 6135
rect 4256 6126 4306 6136
rect 4346 6126 4416 6136
rect 2566 6116 2756 6126
rect 3086 6116 3586 6126
rect 3696 6116 4116 6126
rect 4146 6116 4156 6126
rect 2566 6106 2776 6116
rect 3096 6106 3596 6116
rect 2576 6096 2786 6106
rect 3106 6096 3596 6106
rect 3706 6106 4156 6116
rect 3706 6096 4176 6106
rect 2316 6076 2326 6086
rect 2506 6076 2516 6096
rect 2606 6086 2786 6096
rect 3136 6086 3596 6096
rect 3686 6086 3716 6096
rect 2616 6076 2686 6086
rect 2696 6076 2826 6086
rect 3146 6076 3636 6086
rect 1526 6046 1716 6066
rect 2306 6056 2326 6076
rect 2296 6046 2326 6056
rect 2636 6066 2686 6076
rect 2706 6066 2836 6076
rect 3166 6066 3646 6076
rect 3676 6066 3716 6086
rect 3746 6086 3766 6096
rect 3776 6086 4206 6096
rect 4276 6086 4326 6126
rect 4356 6116 4416 6126
rect 4366 6106 4416 6116
rect 4366 6096 4426 6106
rect 4376 6086 4426 6096
rect 3746 6066 3756 6086
rect 3786 6076 4216 6086
rect 4286 6076 4326 6086
rect 4386 6076 4426 6086
rect 3786 6066 3816 6076
rect 3886 6066 4226 6076
rect 4316 6066 4336 6076
rect 2636 6046 2696 6066
rect 2706 6056 2846 6066
rect 3176 6056 3716 6066
rect 3886 6056 4236 6066
rect 4316 6056 4346 6066
rect 2715 6046 2876 6056
rect 3186 6046 3726 6056
rect 3886 6046 4136 6056
rect 4196 6046 4266 6056
rect 4406 6046 4436 6076
rect 1526 6036 1706 6046
rect 2306 6036 2316 6046
rect 2646 6036 2706 6046
rect 2715 6036 2906 6046
rect 3196 6036 3736 6046
rect 3896 6036 3926 6046
rect 3936 6036 4116 6046
rect 4216 6036 4276 6046
rect 1526 6026 1696 6036
rect 2606 6026 2616 6036
rect 2646 6026 2726 6036
rect 2746 6026 2926 6036
rect 3216 6026 3756 6036
rect 3906 6026 4096 6036
rect 4226 6026 4276 6036
rect 1526 6016 1566 6026
rect 1576 6016 1696 6026
rect 1526 5996 1696 6016
rect 2646 6016 2946 6026
rect 3226 6016 3786 6026
rect 3926 6016 4076 6026
rect 4256 6016 4276 6026
rect 2646 6006 2956 6016
rect 3236 6006 3796 6016
rect 3936 6006 4106 6016
rect 2636 5996 2966 6006
rect 3236 5996 3806 6006
rect 3946 5996 4116 6006
rect 4326 5996 4346 6006
rect 1536 5986 1686 5996
rect 1556 5966 1686 5986
rect 1716 5986 1736 5996
rect 2636 5986 2756 5996
rect 2766 5986 2986 5996
rect 3256 5986 3816 5996
rect 3956 5986 4116 5996
rect 4306 5986 4376 5996
rect 1716 5976 1726 5986
rect 2646 5976 3006 5986
rect 3276 5976 3856 5986
rect 3976 5976 4116 5986
rect 4316 5976 4406 5986
rect 2656 5966 3016 5976
rect 3096 5966 3116 5976
rect 3286 5966 3856 5976
rect 4016 5966 4126 5976
rect 4326 5966 4416 5976
rect 1566 5946 1696 5966
rect 2126 5946 2146 5966
rect 1566 5936 1686 5946
rect 2126 5936 2136 5946
rect 1576 5926 1646 5936
rect 1566 5916 1636 5926
rect 2116 5916 2126 5926
rect 2406 5916 2416 5966
rect 2656 5956 3046 5966
rect 3086 5956 3156 5966
rect 3286 5956 3886 5966
rect 4046 5956 4166 5966
rect 2656 5946 2796 5956
rect 2806 5946 3166 5956
rect 3286 5955 3906 5956
rect 3286 5946 3416 5955
rect 3446 5946 3906 5955
rect 4056 5946 4176 5956
rect 2656 5936 2786 5946
rect 2806 5936 3176 5946
rect 3296 5936 3426 5946
rect 3456 5936 3926 5946
rect 4076 5936 4176 5946
rect 4336 5936 4416 5966
rect 2656 5916 3206 5936
rect 3326 5926 3436 5936
rect 3466 5926 3946 5936
rect 4086 5926 4176 5936
rect 3336 5916 3446 5926
rect 3476 5916 3956 5926
rect 4096 5916 4176 5926
rect 4236 5916 4256 5926
rect 4346 5916 4416 5936
rect 1566 5906 1626 5916
rect 2026 5906 2036 5916
rect 2106 5906 2136 5916
rect 1576 5886 1616 5906
rect 2016 5896 2036 5906
rect 2096 5896 2136 5906
rect 2406 5896 2426 5916
rect 2656 5906 2726 5916
rect 2736 5906 3216 5916
rect 3346 5906 3456 5916
rect 3486 5906 3956 5916
rect 4136 5906 4156 5916
rect 2656 5896 3236 5906
rect 3356 5896 3466 5906
rect 2006 5886 2046 5896
rect 1586 5876 1616 5886
rect 1576 5866 1616 5876
rect 1996 5866 2046 5886
rect 2096 5876 2126 5896
rect 2416 5886 2436 5896
rect 2656 5886 3246 5896
rect 3356 5886 3476 5896
rect 3496 5886 3956 5906
rect 4216 5896 4266 5916
rect 4356 5906 4416 5916
rect 4366 5896 4416 5906
rect 4366 5886 4406 5896
rect 2086 5866 2126 5876
rect 1576 5856 1606 5866
rect 1996 5856 2036 5866
rect 1576 5846 1596 5856
rect 1996 5846 2016 5856
rect 1566 5826 1606 5846
rect 1986 5826 2026 5846
rect 1566 5816 1616 5826
rect 1566 5796 1606 5816
rect 1726 5806 1736 5816
rect 1716 5796 1736 5806
rect 1566 5786 1596 5796
rect 1576 5776 1596 5786
rect 1586 5756 1596 5776
rect 1706 5766 1736 5796
rect 1996 5806 2026 5826
rect 1996 5776 2036 5806
rect 1716 5756 1736 5766
rect 2006 5756 2036 5776
rect 1706 5746 1736 5756
rect 1586 5726 1606 5736
rect 1696 5726 1736 5746
rect 2016 5746 2036 5756
rect 2096 5746 2126 5866
rect 2406 5866 2446 5886
rect 2486 5876 2506 5886
rect 2656 5876 3266 5886
rect 3366 5876 3486 5886
rect 3526 5876 3956 5886
rect 4236 5876 4286 5886
rect 2406 5856 2456 5866
rect 2486 5856 2516 5876
rect 2666 5866 3276 5876
rect 3376 5866 3496 5876
rect 3536 5866 3966 5876
rect 4236 5866 4276 5876
rect 2666 5856 3296 5866
rect 3386 5856 3496 5866
rect 3546 5856 3976 5866
rect 2416 5836 2456 5856
rect 2496 5846 2506 5856
rect 2676 5846 3296 5856
rect 3396 5846 3516 5856
rect 2496 5836 2556 5846
rect 2416 5826 2466 5836
rect 2506 5826 2556 5836
rect 2686 5836 3316 5846
rect 3416 5836 3516 5846
rect 3556 5846 3996 5856
rect 3556 5836 4026 5846
rect 2686 5826 3326 5836
rect 2416 5816 2476 5826
rect 2506 5816 2566 5826
rect 2696 5816 3226 5826
rect 3246 5816 3326 5826
rect 3436 5826 3516 5836
rect 3566 5826 4026 5836
rect 3436 5816 3526 5826
rect 3576 5816 4036 5826
rect 2426 5806 2476 5816
rect 2516 5806 2576 5816
rect 2696 5806 3346 5816
rect 3436 5806 3536 5816
rect 3576 5806 4056 5816
rect 2286 5776 2306 5796
rect 2436 5786 2486 5806
rect 2526 5796 2586 5806
rect 2516 5786 2586 5796
rect 2706 5796 3246 5806
rect 3266 5796 3366 5806
rect 3466 5796 3566 5806
rect 3586 5796 4066 5806
rect 2706 5786 3256 5796
rect 3276 5786 3376 5796
rect 3476 5786 4066 5796
rect 2446 5766 2496 5786
rect 2526 5766 2596 5786
rect 2706 5766 3306 5786
rect 3336 5776 3376 5786
rect 3486 5776 4086 5786
rect 3366 5766 3376 5776
rect 3496 5766 3606 5776
rect 3626 5766 4096 5776
rect 2316 5746 2346 5766
rect 2446 5756 2506 5766
rect 2016 5726 2046 5746
rect 2096 5736 2146 5746
rect 2316 5736 2366 5746
rect 2456 5736 2516 5756
rect 1576 5696 1616 5726
rect 1696 5706 1726 5726
rect 2016 5706 2056 5726
rect 2096 5716 2156 5736
rect 2336 5726 2366 5736
rect 2466 5726 2516 5736
rect 2546 5746 2616 5766
rect 2706 5756 3316 5766
rect 2706 5746 3326 5756
rect 2546 5726 2626 5746
rect 2706 5736 3356 5746
rect 3386 5736 3416 5766
rect 3506 5756 3596 5766
rect 3636 5756 4106 5766
rect 3506 5746 3606 5756
rect 3626 5746 4096 5756
rect 4356 5746 4376 5756
rect 3506 5736 4096 5746
rect 4346 5736 4396 5746
rect 2716 5726 3436 5736
rect 3516 5726 4106 5736
rect 4356 5726 4406 5736
rect 2336 5716 2376 5726
rect 2466 5716 2526 5726
rect 2556 5716 2636 5726
rect 2726 5716 3456 5726
rect 3526 5716 4106 5726
rect 4276 5716 4286 5726
rect 4346 5716 4406 5726
rect 2106 5706 2146 5716
rect 2346 5706 2406 5716
rect 2466 5706 2536 5716
rect 2576 5706 2636 5716
rect 2736 5706 3486 5716
rect 3536 5706 4116 5716
rect 4256 5706 4306 5716
rect 4346 5706 4396 5716
rect 1696 5696 1716 5706
rect 1576 5686 1626 5696
rect 1666 5686 1716 5696
rect 1576 5676 1636 5686
rect 1656 5676 1716 5686
rect 1576 5666 1716 5676
rect 1566 5656 1716 5666
rect 1896 5686 1926 5696
rect 2016 5686 2066 5706
rect 1896 5666 1936 5686
rect 2026 5666 2066 5686
rect 1896 5656 1976 5666
rect 1566 5646 1696 5656
rect 1896 5646 1986 5656
rect 2016 5646 2066 5666
rect 2116 5696 2156 5706
rect 2356 5696 2426 5706
rect 2476 5696 2546 5706
rect 2576 5696 2656 5706
rect 2746 5696 3046 5706
rect 3056 5696 3496 5706
rect 3546 5696 4046 5706
rect 4066 5696 4126 5706
rect 4256 5696 4316 5706
rect 4356 5696 4396 5706
rect 2116 5686 2166 5696
rect 2356 5686 2436 5696
rect 2486 5686 2556 5696
rect 2586 5686 2666 5696
rect 2756 5686 3046 5696
rect 3066 5686 3506 5696
rect 3546 5686 4056 5696
rect 4076 5688 4146 5696
rect 4076 5686 4095 5688
rect 4107 5686 4146 5688
rect 4256 5686 4336 5696
rect 4346 5686 4396 5696
rect 2116 5656 2176 5686
rect 2356 5676 2446 5686
rect 2486 5676 2566 5686
rect 2596 5676 2676 5686
rect 2756 5676 3056 5686
rect 3076 5676 3516 5686
rect 3556 5676 4056 5686
rect 2366 5666 2456 5676
rect 2486 5666 2576 5676
rect 2586 5666 2686 5676
rect 2766 5666 3066 5676
rect 3086 5666 3106 5676
rect 3116 5666 3526 5676
rect 3546 5666 4076 5676
rect 4086 5666 4095 5676
rect 4107 5667 4156 5686
rect 4113 5666 4156 5667
rect 4266 5676 4396 5686
rect 4266 5666 4386 5676
rect 2376 5656 2466 5666
rect 2506 5656 2696 5666
rect 2776 5656 3076 5666
rect 3126 5664 4095 5666
rect 3126 5656 4096 5664
rect 4116 5656 4156 5666
rect 4286 5656 4386 5666
rect 2116 5646 2186 5656
rect 1566 5626 1706 5646
rect 1896 5626 1996 5646
rect 1556 5616 1696 5626
rect 1566 5596 1686 5616
rect 1896 5606 2006 5626
rect 2026 5616 2066 5646
rect 2126 5636 2186 5646
rect 2136 5626 2186 5636
rect 2206 5646 2226 5656
rect 2386 5646 2476 5656
rect 2496 5646 2596 5656
rect 2606 5646 2716 5656
rect 2796 5646 3086 5656
rect 3126 5646 4106 5656
rect 4146 5646 4166 5656
rect 4296 5646 4386 5656
rect 2206 5636 2236 5646
rect 2386 5636 2486 5646
rect 2506 5636 2596 5646
rect 2616 5636 2726 5646
rect 2796 5636 3096 5646
rect 3116 5636 4126 5646
rect 4146 5636 4176 5646
rect 4286 5636 4386 5646
rect 2206 5626 2246 5636
rect 2396 5626 2606 5636
rect 2036 5606 2076 5616
rect 2136 5606 2176 5626
rect 2216 5616 2266 5626
rect 2416 5616 2606 5626
rect 2626 5626 2736 5636
rect 2796 5626 2806 5636
rect 2816 5626 3126 5636
rect 3136 5626 4126 5636
rect 4266 5626 4306 5636
rect 4336 5626 4386 5636
rect 2626 5616 2706 5626
rect 2716 5616 2756 5626
rect 2796 5616 4136 5626
rect 4256 5616 4376 5626
rect 2216 5606 2286 5616
rect 2426 5606 2616 5616
rect 2626 5606 2766 5616
rect 2806 5606 4146 5616
rect 4266 5606 4376 5616
rect 1726 5596 1736 5606
rect 1896 5596 2016 5606
rect 2036 5596 2086 5606
rect 2146 5596 2186 5606
rect 2216 5596 2296 5606
rect 2446 5596 2766 5606
rect 2796 5596 3156 5606
rect 1556 5586 1686 5596
rect 1706 5586 1736 5596
rect 1846 5586 1856 5596
rect 1896 5586 2026 5596
rect 2036 5586 2096 5596
rect 1556 5566 1736 5586
rect 1896 5576 2096 5586
rect 2146 5576 2206 5596
rect 2236 5586 2306 5596
rect 2456 5586 2646 5596
rect 2656 5586 3156 5596
rect 3166 5596 4156 5606
rect 4256 5596 4376 5606
rect 3166 5586 4166 5596
rect 4256 5586 4366 5596
rect 2236 5576 2326 5586
rect 2486 5576 2806 5586
rect 2816 5576 3156 5586
rect 3176 5576 4176 5586
rect 1886 5566 2106 5576
rect 2156 5566 2216 5576
rect 2246 5566 2346 5576
rect 2506 5566 3166 5576
rect 1556 5536 1746 5566
rect 1886 5556 2116 5566
rect 2166 5556 2216 5566
rect 2256 5556 2366 5566
rect 2576 5556 3166 5566
rect 3186 5566 4196 5576
rect 3186 5556 4206 5566
rect 4266 5556 4366 5586
rect 1916 5546 2126 5556
rect 2166 5546 2226 5556
rect 2266 5546 2376 5556
rect 2586 5546 3176 5556
rect 3186 5546 4226 5556
rect 1556 5516 1756 5536
rect 1876 5526 2156 5546
rect 2176 5536 2246 5546
rect 2196 5526 2246 5536
rect 1866 5516 2156 5526
rect 1556 5496 1766 5516
rect 1556 5456 1776 5496
rect 1876 5486 2156 5516
rect 2166 5516 2186 5526
rect 2206 5516 2246 5526
rect 2276 5536 2436 5546
rect 2586 5536 4236 5546
rect 4276 5536 4366 5556
rect 2276 5526 2446 5536
rect 2576 5526 4246 5536
rect 2276 5516 2506 5526
rect 2516 5516 3746 5526
rect 3756 5516 4266 5526
rect 4286 5516 4366 5536
rect 2166 5496 2196 5516
rect 2216 5506 2236 5516
rect 2276 5506 2716 5516
rect 2296 5505 2726 5506
rect 2736 5505 4366 5516
rect 2296 5496 4366 5505
rect 2166 5486 2206 5496
rect 2236 5486 2246 5496
rect 2306 5486 2736 5496
rect 1876 5476 2256 5486
rect 2316 5476 2746 5486
rect 2776 5476 4366 5496
rect 1876 5466 2266 5476
rect 2276 5466 2296 5476
rect 2316 5466 2756 5476
rect 2766 5466 4366 5476
rect 1876 5456 2296 5466
rect 1556 5446 1786 5456
rect 1876 5446 2306 5456
rect 2366 5446 4366 5466
rect 1566 5426 1786 5446
rect 1886 5436 2316 5446
rect 2366 5436 2786 5446
rect 2806 5436 4366 5446
rect 1886 5426 2326 5436
rect 2366 5426 2396 5436
rect 1566 5416 1796 5426
rect 1896 5416 2386 5426
rect 2416 5416 4366 5436
rect 1576 5386 1806 5416
rect 1896 5406 4366 5416
rect 1906 5396 4366 5406
rect 1906 5386 4376 5396
rect 1576 5366 1816 5386
rect 1916 5366 4376 5386
rect 1576 5346 1826 5366
rect 1926 5356 4376 5366
rect 1936 5346 4386 5356
rect 1576 5326 1836 5346
rect 1946 5336 2496 5346
rect 1946 5326 2486 5336
rect 2506 5326 4386 5346
rect 1576 5306 1846 5326
rect 1966 5316 2175 5326
rect 2186 5316 4386 5326
rect 4546 5316 4566 5326
rect 1896 5306 1906 5316
rect 1956 5306 2156 5316
rect 2166 5306 2176 5316
rect 2196 5306 2226 5316
rect 2236 5306 4376 5316
rect 4546 5306 4586 5316
rect 1576 5286 1856 5306
rect 1886 5296 1926 5306
rect 1956 5296 2176 5306
rect 2206 5296 2216 5306
rect 2266 5296 2336 5306
rect 2356 5296 4366 5306
rect 4526 5296 4586 5306
rect 1896 5286 1926 5296
rect 1936 5286 2076 5296
rect 2106 5286 2186 5296
rect 2296 5286 2326 5296
rect 2396 5286 4356 5296
rect 4526 5286 4576 5296
rect 1576 5266 1886 5286
rect 1896 5276 2066 5286
rect 2106 5276 2136 5286
rect 2166 5276 2186 5286
rect 2416 5276 4356 5286
rect 4536 5276 4546 5286
rect 4556 5276 4576 5286
rect 1896 5266 2086 5276
rect 2496 5266 4336 5276
rect 1576 5236 2106 5266
rect 2506 5256 4336 5266
rect 2516 5246 2546 5256
rect 2576 5246 4326 5256
rect 2576 5236 4316 5246
rect 1576 5226 2046 5236
rect 2076 5226 2096 5236
rect 2566 5226 4316 5236
rect 1576 5216 2056 5226
rect 2566 5216 2586 5226
rect 2596 5216 4316 5226
rect 1576 5206 2066 5216
rect 2556 5206 2576 5216
rect 2606 5206 2756 5216
rect 1576 5196 2096 5206
rect 2556 5196 2586 5206
rect 1586 5186 2106 5196
rect 2576 5186 2586 5196
rect 2596 5196 2756 5206
rect 2766 5196 4306 5216
rect 2596 5186 2716 5196
rect 2776 5186 4296 5196
rect 1586 5176 2116 5186
rect 2606 5176 2716 5186
rect 1596 5166 2126 5176
rect 1596 5156 2006 5166
rect 2026 5156 2106 5166
rect 1536 5126 1566 5156
rect 1596 5146 1996 5156
rect 2036 5146 2066 5156
rect 2116 5146 2146 5156
rect 2316 5146 2336 5176
rect 2636 5166 2716 5176
rect 2656 5156 2686 5166
rect 2706 5146 2716 5166
rect 2766 5156 2806 5186
rect 2816 5176 4296 5186
rect 2826 5166 4266 5176
rect 2826 5156 4236 5166
rect 2826 5146 4086 5156
rect 4096 5146 4236 5156
rect 1606 5136 1996 5146
rect 2126 5136 2136 5146
rect 2846 5136 4086 5146
rect 4106 5136 4236 5146
rect 1616 5126 1976 5136
rect 2866 5126 4096 5136
rect 1536 5096 1576 5126
rect 1626 5116 1966 5126
rect 2886 5116 4096 5126
rect 4116 5126 4226 5136
rect 4116 5116 4216 5126
rect 1626 5096 1956 5116
rect 2326 5106 2356 5116
rect 2906 5106 4106 5116
rect 4116 5106 4206 5116
rect 1526 5066 1576 5096
rect 1636 5086 1956 5096
rect 2276 5096 2416 5106
rect 2456 5096 2476 5106
rect 2926 5096 4206 5106
rect 2276 5086 2536 5096
rect 2936 5086 4136 5096
rect 1636 5076 1946 5086
rect 2266 5076 2596 5086
rect 2976 5076 4136 5086
rect 4146 5086 4196 5096
rect 4146 5076 4186 5086
rect 1516 5036 1576 5066
rect 1656 5066 1936 5076
rect 2176 5066 2186 5076
rect 2266 5066 2616 5076
rect 3056 5066 4176 5076
rect 1656 5056 1926 5066
rect 2166 5056 2226 5066
rect 2306 5056 2636 5066
rect 3126 5056 3146 5066
rect 3156 5056 4156 5066
rect 1506 5026 1576 5036
rect 1646 5046 1926 5056
rect 2186 5046 2216 5056
rect 2346 5046 2656 5056
rect 2666 5046 2686 5056
rect 3166 5046 4146 5056
rect 1646 5036 1916 5046
rect 2356 5036 2706 5046
rect 3176 5036 4136 5046
rect 1646 5026 1906 5036
rect 2386 5026 2416 5036
rect 2456 5026 2716 5036
rect 3186 5026 4106 5036
rect 1496 5016 1576 5026
rect 1656 5016 1906 5026
rect 2486 5016 2726 5026
rect 3206 5016 4076 5026
rect 1476 5006 1576 5016
rect 1666 5006 1906 5016
rect 2496 5006 2736 5016
rect 3226 5006 4056 5016
rect 1456 4986 1576 5006
rect 1676 4996 1906 5006
rect 2536 4996 2736 5006
rect 3276 4996 4036 5006
rect 4326 4996 4346 5006
rect 1676 4986 1896 4996
rect 2546 4986 2746 4996
rect 3296 4986 4046 4996
rect 1476 4976 1496 4986
rect 1506 4976 1576 4986
rect 1686 4976 1896 4986
rect 2596 4976 2766 4986
rect 3316 4976 4066 4986
rect 4336 4976 4346 4996
rect 1686 4966 1886 4976
rect 2616 4966 2776 4976
rect 3336 4966 4066 4976
rect 1696 4956 1886 4966
rect 2626 4956 2776 4966
rect 2806 4956 2816 4966
rect 3356 4956 4066 4966
rect 1706 4896 1886 4956
rect 2656 4946 2786 4956
rect 2806 4946 2826 4956
rect 3516 4946 4066 4956
rect 2336 4936 2486 4946
rect 2696 4936 2716 4946
rect 2736 4936 2786 4946
rect 3486 4936 3496 4946
rect 3506 4936 3836 4946
rect 3846 4936 4076 4946
rect 2316 4926 2526 4936
rect 2746 4926 2776 4936
rect 3466 4926 3776 4936
rect 3796 4926 3806 4936
rect 3926 4926 4076 4936
rect 2286 4916 2586 4926
rect 3476 4916 3726 4926
rect 3966 4916 4076 4926
rect 2256 4906 2666 4916
rect 3476 4906 3696 4916
rect 3986 4906 4066 4916
rect 2246 4896 2696 4906
rect 3546 4896 3596 4906
rect 3616 4896 3646 4906
rect 1706 4846 1876 4896
rect 2236 4886 2716 4896
rect 3546 4886 3576 4896
rect 2226 4876 2746 4886
rect 2226 4866 2756 4876
rect 2236 4856 2766 4866
rect 2246 4846 2786 4856
rect 3586 4846 3636 4856
rect 1716 4836 1866 4846
rect 1726 4826 1866 4836
rect 1736 4796 1866 4826
rect 2246 4836 2806 4846
rect 3536 4836 3816 4846
rect 2246 4816 2816 4836
rect 3526 4826 3896 4836
rect 3516 4816 3916 4826
rect 2256 4806 2826 4816
rect 3496 4806 3936 4816
rect 2276 4796 2386 4806
rect 2426 4796 2826 4806
rect 3476 4796 3946 4806
rect 1736 4686 1856 4796
rect 2316 4786 2396 4796
rect 2426 4786 2686 4796
rect 2706 4786 2836 4796
rect 3466 4786 3956 4796
rect 2316 4776 2416 4786
rect 2346 4766 2416 4776
rect 2426 4766 2676 4786
rect 2716 4776 2846 4786
rect 3446 4776 3966 4786
rect 2716 4766 2856 4776
rect 3436 4766 3976 4776
rect 2366 4756 2656 4766
rect 2726 4756 2866 4766
rect 3426 4756 3986 4766
rect 2366 4746 2646 4756
rect 2376 4736 2646 4746
rect 2736 4736 2866 4756
rect 3416 4746 3996 4756
rect 3406 4736 3816 4746
rect 3836 4736 3996 4746
rect 2386 4726 2626 4736
rect 2716 4726 2856 4736
rect 3396 4726 3526 4736
rect 3566 4726 3816 4736
rect 3856 4726 3986 4736
rect 2446 4716 2616 4726
rect 2676 4716 2856 4726
rect 3386 4716 3516 4726
rect 3566 4716 3806 4726
rect 3866 4716 4006 4726
rect 2496 4706 2646 4716
rect 2686 4706 2856 4716
rect 2516 4696 2606 4706
rect 2616 4696 2656 4706
rect 2726 4696 2736 4706
rect 2826 4696 2856 4706
rect 3396 4706 3496 4716
rect 3576 4706 3796 4716
rect 2536 4686 2596 4696
rect 2626 4686 2656 4696
rect 3396 4686 3486 4706
rect 3586 4696 3796 4706
rect 3886 4706 4006 4716
rect 3886 4696 3986 4706
rect 3586 4686 3786 4696
rect 3876 4686 3976 4696
rect 1746 4666 1856 4686
rect 2566 4676 2586 4686
rect 3406 4676 3436 4686
rect 3446 4676 3496 4686
rect 3596 4676 3776 4686
rect 3876 4676 3916 4686
rect 3416 4666 3426 4676
rect 3446 4666 3506 4676
rect 3606 4666 3766 4676
rect 3866 4666 3896 4676
rect 1756 4626 1846 4666
rect 3616 4656 3766 4666
rect 3856 4656 3886 4666
rect 3616 4646 3746 4656
rect 1766 4606 1846 4626
rect 3586 4636 3746 4646
rect 3586 4616 3716 4636
rect 3736 4626 3756 4636
rect 3736 4616 3776 4626
rect 3586 4606 3626 4616
rect 3756 4606 3766 4616
rect 1776 4576 1806 4606
rect 1816 4596 1836 4606
rect 1786 4566 1806 4576
rect 1796 4556 1816 4566
rect 1796 4456 1806 4476
rect 1796 4436 1816 4456
rect 1806 4426 1816 4436
rect 1816 4406 1836 4416
rect 1826 4396 1836 4406
rect 1806 4296 1836 4306
rect 1816 4276 1836 4296
rect 1806 4226 1836 4246
rect 2706 4226 2726 4236
rect 1816 4216 1826 4226
rect 2696 4216 2766 4226
rect 2686 4206 2766 4216
rect 2676 4196 2776 4206
rect 3416 4196 3456 4206
rect 2626 4186 2776 4196
rect 2606 4166 2776 4186
rect 3406 4186 3466 4196
rect 3406 4176 3476 4186
rect 2586 4156 2776 4166
rect 2566 4146 2776 4156
rect 2546 4136 2776 4146
rect 2506 4116 2776 4136
rect 3396 4166 3486 4176
rect 3396 4156 3526 4166
rect 3396 4136 3536 4156
rect 3396 4126 3566 4136
rect 3396 4116 3576 4126
rect 1776 4106 1846 4116
rect 2446 4106 2776 4116
rect 1776 4096 1856 4106
rect 2366 4096 2376 4106
rect 1776 4076 1866 4096
rect 2366 4086 2386 4096
rect 2356 4076 2396 4086
rect 2436 4076 2776 4106
rect 3406 4106 3586 4116
rect 1776 4066 1876 4076
rect 2346 4066 2416 4076
rect 2446 4066 2786 4076
rect 1706 4056 1716 4066
rect 1686 4026 1786 4036
rect 1796 4026 1876 4066
rect 2246 4056 2266 4066
rect 2326 4056 2786 4066
rect 2216 4046 2296 4056
rect 2316 4046 2786 4056
rect 2216 4036 2786 4046
rect 2196 4035 2786 4036
rect 3406 4066 3636 4106
rect 4176 4096 4186 4106
rect 4146 4076 4186 4086
rect 4136 4066 4186 4076
rect 3406 4056 3696 4066
rect 4126 4056 4186 4066
rect 4196 4056 4216 4066
rect 3406 4046 3706 4056
rect 4156 4046 4186 4056
rect 3406 4036 3716 4046
rect 4166 4036 4176 4046
rect 2196 4026 2796 4035
rect 3406 4026 3756 4036
rect 1676 4016 1886 4026
rect 2186 4016 2226 4026
rect 2236 4016 2716 4026
rect 2746 4016 2776 4026
rect 2786 4016 2816 4026
rect 3396 4016 3776 4026
rect 4166 4016 4176 4026
rect 1566 4006 1586 4016
rect 1616 4006 1886 4016
rect 1566 3996 1886 4006
rect 2176 4006 2716 4016
rect 2756 4006 2766 4016
rect 2786 4006 2856 4016
rect 3396 4006 3806 4016
rect 3816 4006 3846 4016
rect 4156 4006 4236 4016
rect 2176 3996 2696 4006
rect 1566 3986 1636 3996
rect 1656 3986 1896 3996
rect 1686 3976 1696 3986
rect 1786 3976 1896 3986
rect 2176 3986 2676 3996
rect 2776 3986 2866 4006
rect 3446 3996 3846 4006
rect 3876 3996 3886 4006
rect 4116 3996 4246 4006
rect 3456 3986 3916 3996
rect 2176 3976 2656 3986
rect 2816 3976 2896 3986
rect 3466 3976 3926 3986
rect 4106 3976 4256 3996
rect 1776 3966 1896 3976
rect 1566 3956 1896 3966
rect 2166 3966 2646 3976
rect 2836 3966 2906 3976
rect 3466 3966 3936 3976
rect 2166 3956 2636 3966
rect 2846 3956 2956 3966
rect 3256 3956 3276 3966
rect 3476 3956 3956 3966
rect 1546 3946 1906 3956
rect 1516 3936 1906 3946
rect 2166 3936 2626 3956
rect 2846 3946 2966 3956
rect 2856 3936 2866 3946
rect 1136 3926 1186 3936
rect 1236 3926 1246 3936
rect 1276 3926 1306 3936
rect 1316 3926 1396 3936
rect 1436 3926 1446 3936
rect 1506 3926 1906 3936
rect 2176 3926 2616 3936
rect 2876 3926 2976 3946
rect 3156 3936 3216 3946
rect 3066 3926 3226 3936
rect 3236 3926 3286 3956
rect 3486 3946 3956 3956
rect 4096 3946 4246 3976
rect 3506 3936 3966 3946
rect 4096 3936 4266 3946
rect 3506 3926 3976 3936
rect 4086 3926 4266 3936
rect 1086 3916 1106 3926
rect 1126 3916 1206 3926
rect 1216 3916 1256 3926
rect 1266 3916 1406 3926
rect 1436 3916 1906 3926
rect 2196 3916 2606 3926
rect 2876 3916 2996 3926
rect 3056 3916 3176 3926
rect 3186 3916 3276 3926
rect 3486 3916 3956 3926
rect 4086 3916 4276 3926
rect 1086 3906 1776 3916
rect 1806 3906 1916 3916
rect 1086 3896 1766 3906
rect 1826 3896 1916 3906
rect 2166 3906 2596 3916
rect 2886 3906 3016 3916
rect 3026 3906 3176 3916
rect 3196 3906 3266 3916
rect 3486 3906 3976 3916
rect 2166 3896 2586 3906
rect 2896 3896 3176 3906
rect 3186 3896 3256 3906
rect 1086 3886 1756 3896
rect 1836 3886 1926 3896
rect 2166 3886 2206 3896
rect 2216 3886 2596 3896
rect 2876 3886 2886 3896
rect 2906 3886 3256 3896
rect 1086 3876 1726 3886
rect 1086 3866 1716 3876
rect 1836 3866 1936 3886
rect 2246 3876 2596 3886
rect 2896 3876 3256 3886
rect 3516 3886 3976 3906
rect 4076 3906 4276 3916
rect 4076 3896 4286 3906
rect 4076 3886 4296 3896
rect 3516 3876 3956 3886
rect 4086 3876 4316 3886
rect 1086 3856 1696 3866
rect 1086 3846 1686 3856
rect 1826 3846 1936 3866
rect 2236 3866 2606 3876
rect 2896 3866 3246 3876
rect 3506 3866 3936 3876
rect 4086 3866 4396 3876
rect 2236 3856 2636 3866
rect 2916 3856 2926 3866
rect 2936 3856 3236 3866
rect 3496 3856 3926 3866
rect 4086 3856 4416 3866
rect 2236 3846 2646 3856
rect 2946 3846 3226 3856
rect 3486 3846 3926 3856
rect 4076 3846 4416 3856
rect 1086 3836 1676 3846
rect 1836 3836 1946 3846
rect 2226 3836 2696 3846
rect 2956 3836 3216 3846
rect 3466 3836 3926 3846
rect 4066 3836 4426 3846
rect 1086 3816 1666 3836
rect 1826 3816 1956 3836
rect 2126 3816 2146 3836
rect 2216 3826 2706 3836
rect 2976 3826 3196 3836
rect 3446 3826 3906 3836
rect 2196 3816 2246 3826
rect 2256 3816 2716 3826
rect 2996 3816 3166 3826
rect 3426 3816 3916 3826
rect 1086 3796 1646 3816
rect 1826 3796 1966 3816
rect 2116 3796 2136 3816
rect 2196 3806 2206 3816
rect 2236 3806 2276 3816
rect 2286 3806 2316 3816
rect 2336 3806 2786 3816
rect 3016 3806 3026 3816
rect 3066 3806 3106 3816
rect 3146 3806 3156 3816
rect 3396 3806 3916 3816
rect 4056 3816 4436 3836
rect 4056 3806 4426 3816
rect 2246 3796 2276 3806
rect 2346 3796 2796 3806
rect 2836 3796 2856 3806
rect 3086 3796 3096 3806
rect 3386 3796 3926 3806
rect 1086 3776 1636 3796
rect 1826 3786 1976 3796
rect 2346 3786 2866 3796
rect 2926 3786 2946 3796
rect 2966 3786 2986 3796
rect 3336 3786 3926 3796
rect 4046 3786 4446 3806
rect 1816 3776 1846 3786
rect 1876 3776 1976 3786
rect 2116 3776 2126 3786
rect 2346 3776 2646 3786
rect 1086 3756 1626 3776
rect 1826 3766 1846 3776
rect 1886 3766 1986 3776
rect 1826 3756 1856 3766
rect 1896 3756 1976 3766
rect 2106 3756 2136 3776
rect 2356 3766 2646 3776
rect 2656 3776 3006 3786
rect 3286 3776 3626 3786
rect 3646 3776 3746 3786
rect 3786 3776 3796 3786
rect 3806 3776 3946 3786
rect 2656 3766 2706 3776
rect 2736 3766 3046 3776
rect 3116 3766 3606 3776
rect 3646 3766 3736 3776
rect 3816 3766 3896 3776
rect 3906 3766 3946 3776
rect 4046 3776 4496 3786
rect 4046 3766 4646 3776
rect 2356 3756 2696 3766
rect 2756 3756 3576 3766
rect 1086 3746 1616 3756
rect 1826 3746 1846 3756
rect 1896 3746 1986 3756
rect 2366 3746 2496 3756
rect 2506 3746 2686 3756
rect 2766 3746 3366 3756
rect 3406 3746 3566 3756
rect 3656 3746 3736 3766
rect 3806 3759 3946 3766
rect 3804 3756 3946 3759
rect 4036 3756 4666 3766
rect 3804 3746 3936 3756
rect 4026 3746 4676 3756
rect 1086 3736 1606 3746
rect 1786 3736 1796 3746
rect 1806 3736 1846 3746
rect 1876 3736 1996 3746
rect 2366 3736 2486 3746
rect 2516 3736 2686 3746
rect 2776 3736 3356 3746
rect 3406 3736 3556 3746
rect 3656 3736 3726 3746
rect 3804 3744 3926 3746
rect 3816 3736 3926 3744
rect 4016 3736 4676 3746
rect 1086 3726 1566 3736
rect 1776 3726 1836 3736
rect 1876 3726 2006 3736
rect 2146 3726 2156 3736
rect 1086 3716 1556 3726
rect 1776 3716 1816 3726
rect 1866 3716 2006 3726
rect 2136 3716 2156 3726
rect 2376 3716 2466 3736
rect 2536 3716 2686 3736
rect 2786 3726 3346 3736
rect 3406 3726 3546 3736
rect 3656 3726 3706 3736
rect 3816 3726 3896 3736
rect 4006 3726 4666 3736
rect 2786 3716 3336 3726
rect 3406 3716 3536 3726
rect 3666 3716 3706 3726
rect 3826 3716 3906 3726
rect 4006 3716 4656 3726
rect 1086 3706 1496 3716
rect 1756 3706 1806 3716
rect 1086 3686 1486 3706
rect 1776 3696 1806 3706
rect 1846 3706 2016 3716
rect 1846 3696 2026 3706
rect 2366 3696 2466 3716
rect 2556 3706 2686 3716
rect 2856 3706 3326 3716
rect 3406 3706 3526 3716
rect 3666 3706 3696 3716
rect 3826 3706 3926 3716
rect 1866 3686 2036 3696
rect 1086 3676 1466 3686
rect 1856 3676 2036 3686
rect 2376 3686 2466 3696
rect 2566 3686 2686 3706
rect 2866 3696 2936 3706
rect 2966 3696 3266 3706
rect 3286 3696 3316 3706
rect 3406 3696 3516 3706
rect 3666 3696 3686 3706
rect 3856 3696 3886 3706
rect 3906 3696 3926 3706
rect 1086 3666 1456 3676
rect 1836 3666 2046 3676
rect 1086 3656 1446 3666
rect 1086 3646 1436 3656
rect 1086 3636 1426 3646
rect 1086 3616 1416 3636
rect 1826 3626 2056 3666
rect 2376 3656 2476 3686
rect 2586 3676 2686 3686
rect 2876 3686 2916 3696
rect 2986 3686 3246 3696
rect 3296 3686 3316 3696
rect 3416 3686 3506 3696
rect 3796 3686 3816 3696
rect 3866 3686 3886 3696
rect 3916 3686 3926 3696
rect 3996 3686 4256 3716
rect 2876 3676 2906 3686
rect 3016 3676 3116 3686
rect 3196 3676 3236 3686
rect 3406 3676 3496 3686
rect 3876 3676 3886 3686
rect 3996 3676 4146 3686
rect 4156 3676 4256 3686
rect 2616 3666 2696 3676
rect 2786 3666 2796 3676
rect 2886 3666 2896 3676
rect 3026 3666 3096 3676
rect 3216 3666 3226 3676
rect 3406 3666 3486 3676
rect 3876 3666 3896 3676
rect 3996 3666 4136 3676
rect 4166 3666 4246 3676
rect 2386 3646 2476 3656
rect 2656 3656 2696 3666
rect 2776 3656 2806 3666
rect 2656 3646 2706 3656
rect 2766 3646 2816 3656
rect 2396 3626 2476 3646
rect 2666 3636 2686 3646
rect 2696 3636 2816 3646
rect 3046 3646 3076 3666
rect 3296 3656 3306 3666
rect 3396 3656 3446 3666
rect 3826 3656 3836 3666
rect 3876 3656 3906 3666
rect 4016 3656 4126 3666
rect 4186 3656 4226 3666
rect 3046 3636 3066 3646
rect 3286 3636 3326 3656
rect 3396 3646 3436 3656
rect 3656 3646 3666 3656
rect 3826 3646 3906 3656
rect 4046 3646 4096 3656
rect 3396 3636 3416 3646
rect 3836 3636 3896 3646
rect 2706 3626 2826 3636
rect 3276 3626 3346 3636
rect 3836 3626 3856 3636
rect 1086 3596 1396 3616
rect 1086 3586 1376 3596
rect 1816 3586 2056 3626
rect 2386 3616 2486 3626
rect 2706 3616 2836 3626
rect 3266 3616 3356 3626
rect 3826 3616 3856 3626
rect 2396 3596 2486 3616
rect 2716 3606 2846 3616
rect 2876 3606 2896 3616
rect 3246 3606 3346 3616
rect 3806 3606 3856 3616
rect 3876 3606 3886 3616
rect 2746 3596 2906 3606
rect 3206 3596 3346 3606
rect 3796 3596 3886 3606
rect 2396 3586 2496 3596
rect 2756 3586 2906 3596
rect 1086 3576 1366 3586
rect 1086 3566 1336 3576
rect 1086 3556 1316 3566
rect 1796 3556 2056 3586
rect 2386 3576 2406 3586
rect 2416 3576 2496 3586
rect 2796 3576 2906 3586
rect 3196 3586 3326 3596
rect 3786 3586 3876 3596
rect 3196 3576 3316 3586
rect 3696 3576 3716 3586
rect 2426 3566 2496 3576
rect 2806 3566 2936 3576
rect 3196 3566 3306 3576
rect 2436 3556 2446 3566
rect 2486 3556 2496 3566
rect 2816 3556 2966 3566
rect 3186 3556 3266 3566
rect 3686 3556 3716 3576
rect 3786 3576 3806 3586
rect 3786 3566 3816 3576
rect 3736 3556 3746 3566
rect 3756 3556 3816 3566
rect 3826 3566 3866 3586
rect 3826 3556 3856 3566
rect 1086 3546 1306 3556
rect 1786 3546 2056 3556
rect 1086 3536 1296 3546
rect 1086 3516 1286 3536
rect 1776 3526 2046 3546
rect 2426 3536 2446 3556
rect 2836 3546 3016 3556
rect 3036 3546 3066 3556
rect 3106 3546 3246 3556
rect 2876 3536 3206 3546
rect 2906 3526 3176 3536
rect 3726 3526 3816 3556
rect 1766 3516 2046 3526
rect 2966 3516 3136 3526
rect 3696 3516 3816 3526
rect 1086 3506 1256 3516
rect 1086 3496 1246 3506
rect 1756 3496 2046 3516
rect 3036 3506 3056 3516
rect 3686 3506 3816 3516
rect 1086 3486 1236 3496
rect 1756 3486 2036 3496
rect 2406 3486 2416 3506
rect 3666 3496 3806 3506
rect 3666 3486 3796 3496
rect 1086 3476 1226 3486
rect 1086 3466 1216 3476
rect 1086 3456 1196 3466
rect 1756 3456 2026 3486
rect 2806 3466 2886 3476
rect 3316 3466 3326 3486
rect 3676 3476 3796 3486
rect 3676 3466 3776 3476
rect 3786 3466 3796 3476
rect 2786 3456 2886 3466
rect 3666 3456 3776 3466
rect 1086 3446 1186 3456
rect 1756 3446 2016 3456
rect 2786 3446 2896 3456
rect 3196 3446 3206 3456
rect 3656 3446 3776 3456
rect 3786 3446 3806 3456
rect 1086 3436 1176 3446
rect 1756 3436 2006 3446
rect 1086 3426 1166 3436
rect 1086 3416 1146 3426
rect 1746 3416 2006 3436
rect 2316 3426 2326 3446
rect 2802 3444 2906 3446
rect 2816 3436 2906 3444
rect 3186 3436 3206 3446
rect 3226 3436 3246 3446
rect 3656 3436 3806 3446
rect 3836 3436 3856 3446
rect 2816 3426 2916 3436
rect 2986 3426 3016 3436
rect 3076 3426 3086 3436
rect 3176 3435 3206 3436
rect 3216 3435 3246 3436
rect 3176 3426 3246 3435
rect 2836 3416 2926 3426
rect 2976 3416 3016 3426
rect 3026 3416 3046 3426
rect 3066 3416 3116 3426
rect 3166 3416 3186 3426
rect 3206 3416 3246 3426
rect 3646 3426 3806 3436
rect 3826 3426 3856 3436
rect 3646 3416 3816 3426
rect 1086 3396 1136 3416
rect 1736 3406 2006 3416
rect 2846 3406 2856 3416
rect 2866 3406 2936 3416
rect 2946 3406 3056 3416
rect 3066 3406 3236 3416
rect 3256 3406 3276 3416
rect 3656 3406 3816 3416
rect 1736 3396 1996 3406
rect 1086 3386 1126 3396
rect 1096 3376 1106 3386
rect 1726 3356 1986 3396
rect 2296 3376 2316 3386
rect 2286 3366 2316 3376
rect 2876 3376 3276 3406
rect 3336 3386 3356 3406
rect 3626 3386 3846 3406
rect 3326 3376 3346 3386
rect 3616 3376 3846 3386
rect 2876 3366 2906 3376
rect 2296 3356 2326 3366
rect 2776 3356 2796 3366
rect 2866 3356 2906 3366
rect 2916 3366 3276 3376
rect 3296 3366 3336 3376
rect 3616 3366 3856 3376
rect 2916 3356 3326 3366
rect 1726 3346 1976 3356
rect 2306 3346 2316 3356
rect 2376 3346 2396 3356
rect 1716 3336 1976 3346
rect 2366 3336 2396 3346
rect 2766 3346 2796 3356
rect 2816 3346 2826 3356
rect 2856 3346 3326 3356
rect 3606 3346 3866 3366
rect 2766 3336 2786 3346
rect 2816 3336 3316 3346
rect 3586 3336 3866 3346
rect 1706 3306 1966 3336
rect 2296 3316 2396 3336
rect 2716 3326 2736 3336
rect 2776 3326 2786 3336
rect 2836 3326 3306 3336
rect 3576 3326 3876 3336
rect 2836 3316 3276 3326
rect 3576 3316 3886 3326
rect 2296 3306 2356 3316
rect 2376 3306 2396 3316
rect 2826 3306 3276 3316
rect 3566 3306 3896 3316
rect 1706 3286 1956 3306
rect 2296 3296 2386 3306
rect 2406 3296 2416 3306
rect 2836 3296 3266 3306
rect 3556 3296 3876 3306
rect 3886 3296 3896 3306
rect 1696 3276 1956 3286
rect 2336 3276 2376 3296
rect 2406 3286 2426 3296
rect 2846 3286 3206 3296
rect 3216 3286 3246 3296
rect 2406 3276 2456 3286
rect 2866 3276 2886 3286
rect 2936 3276 3206 3286
rect 1686 3256 1956 3276
rect 2346 3266 2376 3276
rect 2416 3266 2466 3276
rect 2956 3266 3036 3276
rect 3076 3266 3086 3276
rect 3196 3266 3206 3276
rect 3536 3266 3856 3296
rect 2346 3256 2406 3266
rect 2426 3256 2466 3266
rect 3006 3256 3026 3266
rect 3526 3256 3866 3266
rect 1696 3236 1946 3256
rect 2356 3246 2406 3256
rect 2436 3246 2446 3256
rect 1686 3226 1946 3236
rect 2316 3228 2346 3237
rect 2366 3236 2426 3246
rect 3516 3236 3876 3256
rect 2316 3226 2337 3228
rect 2366 3226 2506 3236
rect 3516 3226 3866 3236
rect 1686 3216 1936 3226
rect 2326 3216 2337 3226
rect 2356 3216 2506 3226
rect 3506 3216 3876 3226
rect 1686 3206 1926 3216
rect 2346 3206 2516 3216
rect 3496 3206 3886 3216
rect 1676 3186 1926 3206
rect 1666 3176 1926 3186
rect 2356 3196 2516 3206
rect 3486 3196 3886 3206
rect 2356 3186 2526 3196
rect 2356 3176 2546 3186
rect 3486 3176 3896 3196
rect 1676 3166 1916 3176
rect 2376 3166 2556 3176
rect 3486 3166 3886 3176
rect 1676 3156 1906 3166
rect 1666 3146 1906 3156
rect 1656 3116 1906 3146
rect 2386 3156 2556 3166
rect 3466 3156 3886 3166
rect 2386 3136 2566 3156
rect 3456 3146 3876 3156
rect 2376 3126 2586 3136
rect 3456 3126 3886 3146
rect 2376 3116 2596 3126
rect 3446 3116 3886 3126
rect 1666 3106 1906 3116
rect 2406 3106 2606 3116
rect 1666 3086 1896 3106
rect 2386 3090 2396 3096
rect 2416 3090 2606 3106
rect 3436 3106 3916 3116
rect 3436 3096 3906 3106
rect 2386 3086 2606 3090
rect 3406 3086 3416 3096
rect 3426 3086 3906 3096
rect 1666 3076 1906 3086
rect 2386 3076 2626 3086
rect 3396 3076 3906 3086
rect 1656 3046 1886 3076
rect 2394 3075 2646 3076
rect 2406 3066 2646 3075
rect 3386 3066 3906 3076
rect 2396 3056 2656 3066
rect 3376 3056 3916 3066
rect 2406 3046 2416 3056
rect 2436 3046 2666 3056
rect 3346 3046 3926 3056
rect 1636 3006 1886 3046
rect 2436 3036 2676 3046
rect 2686 3036 2696 3046
rect 3326 3036 3926 3046
rect 2446 3026 2716 3036
rect 3316 3026 3926 3036
rect 2486 3016 2726 3026
rect 3286 3016 3936 3026
rect 2416 3006 2466 3016
rect 2486 3006 2756 3016
rect 3246 3006 3926 3016
rect 1636 2996 1876 3006
rect 2406 2996 2776 3006
rect 3236 2996 3926 3006
rect 1636 2986 1886 2996
rect 2426 2986 2796 2996
rect 2826 2986 2846 2996
rect 2876 2986 2896 2996
rect 2906 2986 2936 2996
rect 2956 2986 3026 2996
rect 3056 2986 3126 2996
rect 3156 2986 3926 2996
rect 1626 2916 1886 2986
rect 2436 2966 2846 2986
rect 2866 2976 3026 2986
rect 3046 2976 3916 2986
rect 2856 2966 3026 2976
rect 3036 2966 3916 2976
rect 2456 2956 3916 2966
rect 2406 2936 2416 2956
rect 2466 2946 3916 2956
rect 2466 2936 3926 2946
rect 2426 2926 2506 2936
rect 2516 2926 3926 2936
rect 2436 2916 2486 2926
rect 2526 2916 3926 2926
rect 1616 2906 1886 2916
rect 2446 2906 2476 2916
rect 2516 2906 3936 2916
rect 1616 2886 1896 2906
rect 2486 2896 3936 2906
rect 2346 2886 2386 2896
rect 2496 2886 3936 2896
rect 1606 2866 1876 2886
rect 2356 2876 2396 2886
rect 2306 2866 2316 2876
rect 2366 2866 2406 2876
rect 2546 2866 3936 2886
rect 1606 2856 1886 2866
rect 2296 2856 2326 2866
rect 2376 2856 2406 2866
rect 2486 2856 3936 2866
rect 1606 2816 1896 2856
rect 2376 2846 2466 2856
rect 2476 2846 3936 2856
rect 2376 2836 3936 2846
rect 2256 2826 2276 2836
rect 2376 2826 2456 2836
rect 2476 2826 3936 2836
rect 2246 2816 2286 2826
rect 2336 2816 2366 2826
rect 2386 2816 2436 2826
rect 2486 2816 3936 2826
rect 1606 2806 1906 2816
rect 2276 2806 2296 2816
rect 2496 2806 3936 2816
rect 3956 2806 3966 2826
rect 1606 2786 1896 2806
rect 2276 2786 2306 2806
rect 2406 2796 2426 2806
rect 2496 2796 3966 2806
rect 2376 2786 2436 2796
rect 1606 2776 1886 2786
rect 1596 2746 1896 2776
rect 2216 2766 2236 2786
rect 2276 2776 2296 2786
rect 2386 2776 2446 2786
rect 2486 2776 2586 2796
rect 2616 2786 3966 2796
rect 2606 2776 3966 2786
rect 2266 2766 2296 2776
rect 2346 2766 2366 2776
rect 2386 2766 2466 2776
rect 2266 2756 2286 2766
rect 2356 2756 2376 2766
rect 2426 2756 2456 2766
rect 2496 2756 3976 2776
rect 2256 2746 2306 2756
rect 2366 2746 2446 2756
rect 2486 2746 3986 2756
rect 1596 2726 1906 2746
rect 2256 2736 2316 2746
rect 2366 2736 3976 2746
rect 2216 2726 2246 2736
rect 2266 2726 2306 2736
rect 2366 2727 2496 2736
rect 1586 2716 1906 2726
rect 2266 2716 2296 2726
rect 2364 2716 2496 2727
rect 2506 2726 3986 2736
rect 2516 2716 3996 2726
rect 1586 2706 1896 2716
rect 2266 2706 2326 2716
rect 2364 2715 2388 2716
rect 2366 2706 2376 2715
rect 2416 2706 4006 2716
rect 1576 2696 1886 2706
rect 2186 2696 2206 2706
rect 2256 2696 2326 2706
rect 2356 2696 2376 2706
rect 2406 2696 4006 2706
rect 1576 2686 1906 2696
rect 1586 2666 1906 2686
rect 2176 2686 2216 2696
rect 2266 2686 2436 2696
rect 2456 2686 4006 2696
rect 2176 2676 2206 2686
rect 2276 2676 4006 2686
rect 2176 2666 2196 2676
rect 1586 2656 1886 2666
rect 2246 2656 2266 2676
rect 2286 2666 4016 2676
rect 2316 2656 4016 2666
rect 1576 2646 1886 2656
rect 2196 2646 2216 2656
rect 1576 2626 1836 2646
rect 2186 2636 2216 2646
rect 2256 2636 4026 2656
rect 1896 2626 1916 2636
rect 2196 2626 2216 2636
rect 2236 2626 2356 2636
rect 2366 2626 4036 2636
rect 1576 2616 1846 2626
rect 1896 2616 1926 2626
rect 2236 2616 4046 2626
rect 1576 2596 1866 2616
rect 2236 2606 2266 2616
rect 2286 2606 4056 2616
rect 2286 2596 4066 2606
rect 1576 2586 1826 2596
rect 2216 2586 2236 2596
rect 2286 2586 4026 2596
rect 4046 2586 4066 2596
rect 1576 2566 1836 2586
rect 2146 2576 2186 2586
rect 2156 2566 2186 2576
rect 2216 2566 2246 2586
rect 2296 2576 4016 2586
rect 1576 2556 1806 2566
rect 2266 2556 2276 2566
rect 2306 2556 3996 2576
rect 1576 2546 1816 2556
rect 1576 2536 1806 2546
rect 2256 2536 3996 2556
rect 4366 2556 4376 2566
rect 4366 2536 4386 2556
rect 1576 2526 1786 2536
rect 2276 2526 3996 2536
rect 1566 2516 1786 2526
rect 2076 2516 2096 2526
rect 1566 2506 1766 2516
rect 2176 2506 2206 2516
rect 2286 2506 2306 2526
rect 2316 2506 4006 2526
rect 1576 2496 1766 2506
rect 2166 2496 2216 2506
rect 1576 2476 1776 2496
rect 2186 2486 2216 2496
rect 2246 2486 2276 2506
rect 2286 2486 4006 2506
rect 2076 2476 2096 2486
rect 2196 2476 2206 2486
rect 1576 2466 1766 2476
rect 1576 2446 1756 2466
rect 2196 2456 2206 2466
rect 2296 2456 2326 2486
rect 2346 2476 4016 2486
rect 4286 2476 4296 2486
rect 4376 2476 4396 2486
rect 2336 2456 4026 2476
rect 4286 2466 4316 2476
rect 4366 2466 4446 2476
rect 4276 2456 4326 2466
rect 4356 2456 4446 2466
rect 2186 2446 2216 2456
rect 2246 2446 2266 2456
rect 2296 2446 4036 2456
rect 4256 2446 4436 2456
rect 1576 2426 1736 2446
rect 2246 2436 2276 2446
rect 2306 2436 2326 2446
rect 2336 2436 2356 2446
rect 2256 2426 2276 2436
rect 2376 2426 4036 2446
rect 4246 2436 4346 2446
rect 4366 2436 4396 2446
rect 4406 2436 4436 2446
rect 4246 2426 4336 2436
rect 4416 2426 4436 2436
rect 1576 2416 1716 2426
rect 2336 2416 2346 2426
rect 2386 2416 4046 2426
rect 4256 2416 4366 2426
rect 1576 2406 1706 2416
rect 2266 2406 2286 2416
rect 1576 2386 1696 2406
rect 2276 2396 2286 2406
rect 2306 2406 4046 2416
rect 4266 2406 4386 2416
rect 2306 2396 2376 2406
rect 1716 2386 1726 2396
rect 2326 2386 2376 2396
rect 2406 2396 4056 2406
rect 4276 2396 4406 2406
rect 4416 2396 4446 2406
rect 2406 2386 2466 2396
rect 2476 2386 4056 2396
rect 4286 2386 4446 2396
rect 1576 2376 1726 2386
rect 2286 2376 2306 2386
rect 2416 2376 2456 2386
rect 2506 2376 4056 2386
rect 4316 2376 4476 2386
rect 1576 2356 1696 2376
rect 2326 2366 2346 2376
rect 1566 2346 1696 2356
rect 2316 2346 2356 2366
rect 2406 2356 2466 2376
rect 2486 2366 4066 2376
rect 4346 2366 4476 2376
rect 2486 2356 2516 2366
rect 2546 2356 2586 2366
rect 2406 2346 2456 2356
rect 2496 2346 2516 2356
rect 2556 2346 2586 2356
rect 2596 2356 4066 2366
rect 4366 2356 4506 2366
rect 2596 2346 4076 2356
rect 4376 2346 4536 2356
rect 1566 2326 1686 2346
rect 2326 2336 2346 2346
rect 2336 2326 2346 2336
rect 2416 2326 2446 2346
rect 2536 2336 3296 2346
rect 3306 2336 4076 2346
rect 4406 2336 4536 2346
rect 2536 2326 2606 2336
rect 2626 2326 3296 2336
rect 3316 2326 4076 2336
rect 4416 2326 4546 2336
rect 1086 2316 1106 2326
rect 1566 2316 1676 2326
rect 2406 2316 2446 2326
rect 2547 2325 2598 2326
rect 1086 2286 1126 2316
rect 1566 2296 1686 2316
rect 2416 2306 2436 2316
rect 2556 2306 2586 2325
rect 2626 2316 4076 2326
rect 4456 2316 4546 2326
rect 2606 2306 3326 2316
rect 3336 2306 4086 2316
rect 4466 2306 4556 2316
rect 4586 2306 4606 2316
rect 2596 2296 2636 2306
rect 2696 2296 2736 2306
rect 2746 2296 3156 2306
rect 1096 2276 1126 2286
rect 1576 2276 1676 2296
rect 2596 2286 2626 2296
rect 2706 2286 2736 2296
rect 2766 2286 2786 2296
rect 2806 2286 2886 2296
rect 2906 2286 3086 2296
rect 3106 2286 3156 2296
rect 3186 2296 4086 2306
rect 4506 2296 4616 2306
rect 3186 2286 3226 2296
rect 3236 2295 4096 2296
rect 2466 2276 2486 2286
rect 2516 2276 2536 2286
rect 2656 2276 2686 2286
rect 2816 2276 2866 2286
rect 2916 2276 3225 2286
rect 3236 2276 3256 2295
rect 3266 2286 4096 2295
rect 4516 2286 4616 2296
rect 3296 2276 4106 2286
rect 4526 2276 4616 2286
rect 1566 2256 1666 2276
rect 2456 2266 2486 2276
rect 2506 2266 2536 2276
rect 2556 2266 2566 2276
rect 2606 2266 2666 2276
rect 2836 2266 2856 2276
rect 2956 2266 3006 2276
rect 2516 2256 2526 2266
rect 2606 2256 2646 2266
rect 2966 2256 3006 2266
rect 3046 2266 3108 2276
rect 3156 2274 3266 2276
rect 3156 2266 3206 2274
rect 3046 2256 3116 2266
rect 3166 2256 3196 2266
rect 3216 2256 3266 2274
rect 3316 2266 4106 2276
rect 4546 2266 4606 2276
rect 1556 2226 1666 2256
rect 2486 2246 2496 2256
rect 2486 2236 2506 2246
rect 2976 2236 3006 2256
rect 3096 2246 3116 2256
rect 3316 2246 4116 2266
rect 4576 2256 4606 2266
rect 2486 2226 2526 2236
rect 1566 2206 1676 2226
rect 2926 2216 2936 2236
rect 2986 2226 3006 2236
rect 3036 2236 3056 2246
rect 3306 2236 4126 2246
rect 3036 2226 3046 2236
rect 3296 2216 4126 2236
rect 3106 2206 3146 2216
rect 3296 2206 4136 2216
rect 1576 2186 1686 2206
rect 3066 2196 3076 2206
rect 3316 2196 4136 2206
rect 3316 2186 4146 2196
rect 1586 2176 1676 2186
rect 3276 2176 4146 2186
rect 1576 2166 1676 2176
rect 3266 2166 4156 2176
rect 1566 2156 1686 2166
rect 1576 2116 1686 2156
rect 3276 2136 4156 2166
rect 1696 2116 1716 2126
rect 1576 2066 1716 2116
rect 3276 2096 4176 2136
rect 3266 2086 4186 2096
rect 3266 2076 4196 2086
rect 1576 2046 1726 2066
rect 3256 2046 4196 2076
rect 1586 2026 1726 2046
rect 3236 2026 4196 2046
rect 1576 2006 1726 2026
rect 3226 2016 4206 2026
rect 3226 2006 4216 2016
rect 1586 1976 1736 2006
rect 3236 1986 4216 2006
rect 3246 1976 4226 1986
rect 1576 1956 1736 1976
rect 3226 1966 4226 1976
rect 1576 1946 1726 1956
rect 3206 1946 4226 1966
rect 1576 1936 1716 1946
rect 3196 1936 4236 1946
rect 1566 1916 1716 1936
rect 3186 1926 4236 1936
rect 3186 1916 4246 1926
rect 1556 1886 1716 1916
rect 3196 1906 4246 1916
rect 1546 1866 1716 1886
rect 3186 1896 4246 1906
rect 3186 1876 4256 1896
rect 1536 1856 1716 1866
rect 3176 1866 4256 1876
rect 1526 1846 1706 1856
rect 3176 1846 4266 1866
rect 1466 1836 1486 1846
rect 1456 1806 1496 1836
rect 1366 1786 1396 1806
rect 1446 1796 1486 1806
rect 1436 1786 1476 1796
rect 1426 1776 1466 1786
rect 1416 1766 1466 1776
rect 1416 1756 1456 1766
rect 1406 1746 1446 1756
rect 1396 1736 1436 1746
rect 1316 1726 1346 1736
rect 1306 1706 1346 1726
rect 1386 1726 1426 1736
rect 1386 1716 1416 1726
rect 1386 1706 1396 1716
rect 1306 1696 1356 1706
rect 1526 1696 1686 1846
rect 3176 1836 4276 1846
rect 3166 1806 4276 1836
rect 3156 1786 4286 1806
rect 3126 1776 4296 1786
rect 3116 1756 4296 1776
rect 3106 1736 4296 1756
rect 3106 1716 4306 1736
rect 3096 1706 4316 1716
rect 3076 1696 4316 1706
rect 1306 1686 1336 1696
rect 1286 1666 1336 1686
rect 1276 1656 1336 1666
rect 1526 1656 1666 1696
rect 3066 1686 4326 1696
rect 3056 1676 4326 1686
rect 3046 1656 4326 1676
rect 1266 1636 1286 1656
rect 1306 1646 1336 1656
rect 1306 1636 1326 1646
rect 1276 1626 1316 1636
rect 1216 1616 1246 1626
rect 1276 1616 1306 1626
rect 1206 1606 1246 1616
rect 1516 1606 1666 1656
rect 3036 1636 4336 1656
rect 3026 1626 4346 1636
rect 3006 1606 4346 1626
rect 1196 1596 1276 1606
rect 1196 1586 1266 1596
rect 1196 1576 1256 1586
rect 1516 1576 1656 1606
rect 3006 1586 4356 1606
rect 2986 1576 4356 1586
rect 1206 1566 1236 1576
rect 1516 1566 1666 1576
rect 2976 1566 4366 1576
rect 1206 1556 1226 1566
rect 1126 1546 1136 1556
rect 1166 1546 1176 1556
rect 1116 1536 1146 1546
rect 1106 1526 1146 1536
rect 1516 1536 1676 1566
rect 2966 1556 4366 1566
rect 2946 1546 4366 1556
rect 2926 1536 4376 1546
rect 1516 1516 1686 1536
rect 2926 1526 4386 1536
rect 1506 1476 1686 1516
rect 2946 1506 4386 1526
rect 2926 1486 4396 1506
rect 2896 1476 4396 1486
rect 1506 1466 1696 1476
rect 1506 1446 1706 1466
rect 2886 1456 4406 1476
rect 1506 1386 1716 1446
rect 2886 1436 4416 1456
rect 2856 1426 4416 1436
rect 2826 1416 4416 1426
rect 2826 1406 4426 1416
rect 2836 1386 4426 1406
rect 1506 1376 1756 1386
rect 2826 1376 4436 1386
rect 1506 1356 1746 1376
rect 2826 1366 4446 1376
rect 1506 1346 1756 1356
rect 2816 1346 4446 1366
rect 1506 1336 1766 1346
rect 2806 1336 4446 1346
rect 1506 1306 1776 1336
rect 2796 1326 4456 1336
rect 2786 1316 4456 1326
rect 1506 1296 1766 1306
rect 2776 1296 4466 1316
rect 1506 1286 1776 1296
rect 2766 1286 4476 1296
rect 1506 1266 1786 1286
rect 2706 1266 2726 1276
rect 2746 1266 4476 1286
rect 1516 1257 1826 1266
rect 1516 1246 1845 1257
rect 2696 1256 4486 1266
rect 2686 1246 4486 1256
rect 1516 1245 1856 1246
rect 1516 1236 1816 1245
rect 1836 1236 1856 1245
rect 2666 1236 4486 1246
rect 1506 1226 1856 1236
rect 2656 1226 4476 1236
rect 1506 1216 1836 1226
rect 2646 1216 4466 1226
rect 1516 1186 1836 1216
rect 2636 1206 4466 1216
rect 2616 1196 4456 1206
rect 2606 1186 4456 1196
rect 1516 1176 1866 1186
rect 2606 1176 4446 1186
rect 1516 1166 1886 1176
rect 1516 1136 1906 1166
rect 2596 1156 4446 1176
rect 2586 1146 4436 1156
rect 2566 1136 4446 1146
rect 1516 1126 1896 1136
rect 2546 1126 4446 1136
rect 1516 1116 1916 1126
rect 2536 1116 4446 1126
rect 1516 1086 1936 1116
rect 2526 1106 4456 1116
rect 2496 1096 4456 1106
rect 1986 1086 1996 1096
rect 2486 1086 4466 1096
rect 1506 1076 1946 1086
rect 2486 1076 4476 1086
rect 1506 1066 1956 1076
rect 2476 1066 4476 1076
rect 1506 1056 1976 1066
rect 2436 1056 4476 1066
rect 1506 1046 2006 1056
rect 2426 1046 4476 1056
rect 1506 1036 2026 1046
rect 2286 1036 2316 1046
rect 2366 1036 4476 1046
rect 1506 1026 2056 1036
rect 1506 1016 2086 1026
rect 2206 1016 2236 1026
rect 2266 1016 2326 1036
rect 2356 1026 4486 1036
rect 2346 1016 4496 1026
rect 1506 1006 2126 1016
rect 2206 1006 2246 1016
rect 2256 1006 4496 1016
rect 1506 996 2136 1006
rect 2216 996 4496 1006
rect 1506 976 4486 996
rect 1506 956 4516 976
rect 1506 946 4526 956
rect 1506 906 4536 946
rect 1506 876 4546 906
rect 1506 866 4556 876
rect 1496 846 4566 866
rect 1496 826 4576 846
rect 1496 786 4586 826
rect 1496 763 4596 786
<< end >>
