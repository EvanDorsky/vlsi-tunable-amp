magic
tech scmos
timestamp 1418768571
<< nwell >>
rect 58 0 62 3
rect 43 -4 86 0
rect 142 0 146 1
rect 129 -4 172 0
rect 0 -136 2 -4
rect 58 -5 62 -4
rect 153 -5 157 -4
<< pwell >>
rect 0 -4 43 3
rect 86 -4 129 3
rect 0 -388 2 -136
<< pdcontact >>
rect 11 -14 15 -10
rect 103 -14 107 -10
<< polysilicon >>
rect 57 3 63 4
rect 109 3 115 4
<< polycontact >>
rect 26 1 30 5
rect 58 -1 62 3
rect 110 -1 114 3
rect 142 1 146 5
rect 153 -9 157 -5
<< metal1 >>
rect 26 -1 30 1
rect 11 -5 30 -1
rect 58 -5 62 -1
rect 103 -5 114 -1
rect 142 0 146 1
rect 142 -4 157 0
rect 153 -5 157 -4
rect 11 -10 15 -5
rect 103 -10 107 -5
use amp  amp_0
timestamp 1418768421
transform 1 0 95 0 1 135
box -95 -135 77 126
use bias  bias_0
timestamp 1418768461
transform 1 0 -11 0 1 -106
box 13 -282 183 102
<< end >>
