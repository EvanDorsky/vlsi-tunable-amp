magic
tech scmos
magscale 1 3
timestamp 1419145638
<< error_p >>
rect 3429 3917 3430 3927
rect 3429 3797 3430 3826
<< metal1 >>
rect 1811 7437 1841 7457
rect 1801 7427 1841 7437
rect 1921 7427 1931 7437
rect 1801 7417 1831 7427
rect 1871 7417 1881 7427
rect 1641 7407 1651 7417
rect 1631 7397 1651 7407
rect 1941 7397 1961 7407
rect 1341 7387 1351 7397
rect 1501 7387 1521 7397
rect 1621 7387 1651 7397
rect 1911 7387 1971 7397
rect 1981 7387 2001 7397
rect 2041 7387 2061 7397
rect 1491 7377 1521 7387
rect 1901 7377 1961 7387
rect 1981 7377 2011 7387
rect 2021 7377 2071 7387
rect 1111 7367 1141 7377
rect 1331 7367 1341 7377
rect 1471 7367 1511 7377
rect 1891 7367 1951 7377
rect 1081 7357 1091 7367
rect 1111 7347 1131 7367
rect 1481 7357 1501 7367
rect 1881 7357 1951 7367
rect 1981 7367 2101 7377
rect 2161 7367 2171 7377
rect 1981 7357 2141 7367
rect 1481 7347 1491 7357
rect 1591 7347 1631 7357
rect 1671 7347 1711 7357
rect 1861 7347 1921 7357
rect 1031 7317 1041 7337
rect 1091 7307 1131 7347
rect 1431 7337 1451 7347
rect 1581 7337 1631 7347
rect 1661 7337 1711 7347
rect 1851 7337 1901 7347
rect 1941 7337 2171 7357
rect 1421 7327 1451 7337
rect 1521 7327 1531 7337
rect 1561 7327 1611 7337
rect 1411 7317 1441 7327
rect 1551 7326 1611 7327
rect 1651 7327 1701 7337
rect 1831 7327 1871 7337
rect 1921 7327 2181 7337
rect 1551 7317 1602 7326
rect 1651 7317 1681 7327
rect 1821 7317 1861 7327
rect 1911 7317 2181 7327
rect 1391 7307 1421 7317
rect 1521 7307 1581 7317
rect 1611 7307 1621 7317
rect 1641 7307 1671 7317
rect 1811 7307 1841 7317
rect 1901 7307 2071 7317
rect 2091 7307 2111 7317
rect 2121 7307 2191 7317
rect 2301 7307 2331 7317
rect 1091 7287 1121 7307
rect 1081 7267 1121 7287
rect 1321 7287 1341 7307
rect 1391 7297 1401 7307
rect 1461 7297 1481 7307
rect 1511 7297 1571 7307
rect 1611 7297 1671 7307
rect 1801 7297 1831 7307
rect 1881 7297 1971 7307
rect 1991 7297 2011 7307
rect 2121 7297 2141 7307
rect 2151 7297 2211 7307
rect 2261 7297 2331 7307
rect 1371 7287 1381 7297
rect 1451 7287 1561 7297
rect 1601 7287 1661 7297
rect 1801 7287 1821 7297
rect 1871 7287 1941 7297
rect 2131 7287 2141 7297
rect 2161 7287 2171 7297
rect 2231 7287 2331 7297
rect 1321 7277 1331 7287
rect 1361 7277 1381 7287
rect 1431 7277 1561 7287
rect 1571 7277 1651 7287
rect 1851 7277 1921 7287
rect 2091 7277 2101 7287
rect 2221 7277 2361 7287
rect 1291 7267 1331 7277
rect 1351 7267 1371 7277
rect 1071 7257 1111 7267
rect 1281 7257 1371 7267
rect 1421 7267 1601 7277
rect 1841 7267 1881 7277
rect 1991 7267 2011 7277
rect 2081 7267 2111 7277
rect 1421 7257 1591 7267
rect 1651 7257 1671 7267
rect 1731 7257 1751 7267
rect 1821 7257 1861 7267
rect 1981 7257 2001 7267
rect 2071 7257 2111 7267
rect 1071 7247 1091 7257
rect 1271 7247 1361 7257
rect 991 7237 1001 7247
rect 1061 7227 1091 7247
rect 1261 7237 1361 7247
rect 1411 7247 1591 7257
rect 1631 7247 1641 7257
rect 1721 7247 1741 7257
rect 1811 7247 1841 7257
rect 1961 7247 2001 7257
rect 2031 7247 2061 7257
rect 2091 7247 2101 7257
rect 2131 7247 2151 7277
rect 2221 7267 2241 7277
rect 2251 7275 2271 7277
rect 2211 7266 2241 7267
rect 2262 7267 2271 7275
rect 2281 7267 2301 7277
rect 2262 7266 2301 7267
rect 2211 7257 2251 7266
rect 2261 7257 2301 7266
rect 2321 7266 2371 7277
rect 2321 7257 2358 7266
rect 2191 7247 2311 7257
rect 2331 7247 2358 7257
rect 1411 7245 1581 7247
rect 1411 7237 1569 7245
rect 1601 7237 1641 7247
rect 1701 7237 1731 7247
rect 1801 7237 1831 7247
rect 1961 7237 2051 7247
rect 2191 7237 2321 7247
rect 2391 7245 2401 7247
rect 2371 7237 2401 7245
rect 1231 7227 1351 7237
rect 1411 7227 1551 7237
rect 1590 7236 1651 7237
rect 1581 7227 1651 7236
rect 1691 7227 1731 7237
rect 1791 7227 1811 7237
rect 1921 7227 1931 7237
rect 1941 7227 2001 7237
rect 2011 7227 2021 7237
rect 2081 7227 2111 7237
rect 2181 7227 2331 7237
rect 2361 7227 2441 7237
rect 881 7217 891 7227
rect 1061 7217 1081 7227
rect 1221 7217 1341 7227
rect 1391 7217 1551 7227
rect 851 7207 901 7217
rect 831 7197 901 7207
rect 811 7177 901 7197
rect 1051 7187 1071 7217
rect 1221 7207 1331 7217
rect 1371 7207 1541 7217
rect 1571 7207 1631 7227
rect 1681 7217 1722 7227
rect 1671 7207 1722 7217
rect 1761 7207 1771 7227
rect 1911 7217 1991 7227
rect 2071 7217 2121 7227
rect 2181 7217 2351 7227
rect 2371 7217 2431 7227
rect 2491 7217 2511 7227
rect 1851 7207 1881 7217
rect 1901 7207 1971 7217
rect 2041 7207 2051 7217
rect 2061 7207 2121 7217
rect 1221 7187 1321 7207
rect 1361 7197 1539 7207
rect 1561 7197 1591 7207
rect 1601 7197 1631 7207
rect 1651 7197 1722 7207
rect 1731 7206 1743 7207
rect 1731 7197 1751 7206
rect 1801 7197 1811 7207
rect 1851 7197 1871 7207
rect 1891 7197 1931 7207
rect 2041 7197 2111 7207
rect 1351 7187 1539 7197
rect 1551 7187 1581 7197
rect 1041 7177 1071 7187
rect 1211 7177 1311 7187
rect 1341 7177 1591 7187
rect 1601 7177 1691 7197
rect 1711 7187 1751 7197
rect 1841 7187 1861 7197
rect 1891 7187 1921 7197
rect 2031 7187 2111 7197
rect 2171 7197 2211 7217
rect 2231 7207 2361 7217
rect 2371 7207 2421 7217
rect 2231 7197 2401 7207
rect 2481 7197 2502 7217
rect 2171 7187 2261 7197
rect 2281 7187 2391 7197
rect 2441 7187 2471 7197
rect 2491 7187 2501 7197
rect 2511 7187 2531 7197
rect 2571 7187 2581 7197
rect 1721 7179 1751 7187
rect 1721 7177 1749 7179
rect 801 7167 891 7177
rect 921 7167 931 7177
rect 811 7157 901 7167
rect 921 7157 941 7167
rect 1041 7157 1061 7177
rect 1171 7167 1321 7177
rect 1331 7167 1681 7177
rect 1711 7167 1741 7177
rect 1821 7167 1851 7187
rect 2011 7177 2111 7187
rect 2161 7177 2241 7187
rect 2281 7177 2401 7187
rect 2411 7177 2481 7187
rect 1991 7176 2111 7177
rect 1991 7167 2100 7176
rect 2281 7167 2471 7177
rect 1161 7157 1681 7167
rect 1710 7158 1741 7167
rect 1731 7157 1741 7158
rect 1811 7157 1841 7167
rect 1971 7157 2001 7167
rect 2011 7157 2081 7167
rect 811 7137 891 7157
rect 781 7127 891 7137
rect 911 7137 931 7157
rect 1031 7147 1061 7157
rect 1091 7147 1101 7157
rect 1031 7137 1051 7147
rect 911 7127 941 7137
rect 761 7097 881 7127
rect 901 7107 941 7127
rect 991 7107 1001 7117
rect 891 7097 941 7107
rect 981 7098 1001 7107
rect 1021 7097 1051 7137
rect 1081 7117 1101 7147
rect 771 7077 941 7097
rect 1011 7086 1051 7097
rect 1071 7087 1101 7117
rect 1161 7147 1671 7157
rect 1161 7117 1291 7147
rect 1311 7137 1671 7147
rect 1731 7155 1749 7157
rect 1731 7146 1761 7155
rect 1811 7147 1831 7157
rect 1921 7147 1991 7157
rect 1721 7137 1761 7146
rect 1801 7137 1821 7147
rect 1911 7137 1951 7147
rect 1971 7137 1981 7147
rect 2021 7137 2081 7157
rect 2111 7157 2121 7167
rect 2131 7157 2161 7167
rect 2281 7157 2301 7167
rect 2111 7147 2141 7157
rect 2201 7147 2211 7157
rect 2291 7147 2301 7157
rect 2101 7137 2131 7147
rect 2191 7137 2221 7147
rect 2281 7137 2301 7147
rect 2322 7157 2331 7167
rect 2341 7157 2391 7167
rect 2322 7147 2371 7157
rect 2511 7147 2561 7157
rect 2322 7137 2331 7147
rect 2491 7137 2601 7147
rect 1311 7127 1601 7137
rect 1611 7128 1661 7137
rect 1611 7127 1674 7128
rect 1691 7127 1701 7137
rect 1721 7127 1751 7137
rect 1301 7117 1731 7127
rect 1841 7117 1851 7137
rect 1911 7127 1941 7137
rect 2011 7127 2071 7137
rect 1161 7097 1731 7117
rect 1781 7107 1791 7117
rect 1821 7107 1851 7117
rect 2001 7117 2061 7127
rect 2091 7117 2121 7137
rect 2181 7127 2211 7137
rect 2271 7127 2301 7137
rect 2471 7127 2611 7137
rect 2181 7117 2201 7127
rect 2271 7117 2281 7127
rect 2441 7117 2621 7127
rect 2001 7107 2051 7117
rect 2091 7107 2111 7117
rect 2171 7107 2191 7117
rect 2241 7107 2251 7117
rect 2401 7107 2631 7117
rect 1811 7097 1841 7107
rect 1991 7097 2051 7107
rect 2081 7097 2111 7107
rect 2401 7097 2531 7107
rect 2551 7097 2661 7107
rect 1151 7087 1731 7097
rect 1771 7087 1781 7097
rect 1001 7077 1051 7086
rect 761 7067 951 7077
rect 981 7067 1051 7077
rect 1061 7067 1101 7087
rect 1141 7077 1701 7087
rect 1710 7086 1731 7087
rect 1721 7077 1731 7086
rect 1761 7077 1781 7087
rect 1801 7087 1841 7097
rect 1801 7077 1821 7087
rect 1981 7077 2041 7097
rect 2081 7077 2101 7097
rect 2391 7087 2451 7097
rect 2381 7080 2441 7087
rect 2469 7086 2521 7097
rect 2551 7087 2671 7097
rect 2370 7077 2441 7080
rect 2471 7077 2521 7086
rect 2541 7077 2681 7087
rect 1131 7067 1731 7077
rect 1751 7067 1811 7077
rect 1971 7067 2031 7077
rect 2370 7067 2411 7077
rect 2471 7067 2511 7077
rect 2541 7067 2691 7077
rect 771 6997 951 7067
rect 971 7047 991 7067
rect 1001 7037 1041 7067
rect 1061 7057 1701 7067
rect 1061 7047 1681 7057
rect 1691 7047 1701 7057
rect 991 7027 1041 7037
rect 1051 7037 1701 7047
rect 1721 7047 1831 7067
rect 1971 7057 2021 7067
rect 2370 7065 2394 7067
rect 2370 7057 2381 7065
rect 2471 7062 2501 7067
rect 2001 7047 2011 7057
rect 2081 7047 2091 7057
rect 2361 7050 2381 7057
rect 1721 7037 1821 7047
rect 1991 7037 2011 7047
rect 2071 7037 2091 7047
rect 2346 7047 2381 7050
rect 2460 7047 2501 7062
rect 2541 7057 2701 7067
rect 2531 7047 2691 7057
rect 2346 7037 2371 7047
rect 2441 7037 2471 7047
rect 2481 7037 2491 7047
rect 2521 7037 2641 7047
rect 2661 7037 2681 7047
rect 1051 7027 1791 7037
rect 1981 7027 2001 7037
rect 2061 7027 2081 7037
rect 2341 7035 2370 7037
rect 2341 7027 2361 7035
rect 2431 7027 2471 7037
rect 2521 7027 2631 7037
rect 991 7007 1771 7027
rect 1891 7007 1901 7017
rect 1961 7007 1991 7027
rect 2061 7017 2071 7027
rect 2331 7017 2351 7027
rect 2431 7017 2451 7027
rect 2501 7017 2661 7027
rect 2331 7007 2341 7017
rect 2411 7007 2441 7017
rect 2501 7007 2521 7017
rect 2551 7007 2601 7017
rect 2621 7007 2651 7017
rect 2751 7007 2781 7017
rect 991 6997 1761 7007
rect 1851 6997 1861 7007
rect 1881 6997 1901 7007
rect 1951 6997 1981 7007
rect 2391 6997 2421 7007
rect 751 6977 961 6997
rect 991 6977 1751 6997
rect 1791 6987 1801 6997
rect 1841 6996 1861 6997
rect 1871 6996 1891 6997
rect 1841 6987 1891 6996
rect 1951 6987 1971 6997
rect 2381 6987 2421 6997
rect 2561 6997 2601 7007
rect 2631 6997 2651 7007
rect 2731 6997 2781 7007
rect 2561 6987 2591 6997
rect 2721 6987 2771 6997
rect 1771 6977 1801 6987
rect 761 6967 961 6977
rect 771 6947 961 6967
rect 761 6937 961 6947
rect 751 6927 961 6937
rect 981 6957 1741 6977
rect 1761 6967 1801 6977
rect 1848 6972 1881 6987
rect 2371 6977 2421 6987
rect 2461 6977 2481 6987
rect 2511 6977 2571 6987
rect 2711 6977 2751 6987
rect 1851 6967 1881 6972
rect 2051 6967 2071 6977
rect 2301 6967 2331 6977
rect 2361 6967 2412 6977
rect 1751 6957 1791 6967
rect 1851 6957 1871 6967
rect 1941 6957 1981 6967
rect 2031 6957 2071 6967
rect 2291 6957 2321 6967
rect 2351 6966 2412 6967
rect 2451 6967 2481 6977
rect 2501 6967 2561 6977
rect 2691 6967 2731 6977
rect 2351 6957 2381 6966
rect 981 6947 1041 6957
rect 1051 6947 1791 6957
rect 1841 6947 1871 6957
rect 1921 6947 1981 6957
rect 2011 6947 2061 6957
rect 2281 6947 2311 6957
rect 2341 6947 2371 6957
rect 2401 6947 2411 6966
rect 2451 6957 2561 6967
rect 2671 6957 2721 6967
rect 2451 6947 2511 6957
rect 2541 6947 2561 6957
rect 2661 6947 2701 6957
rect 981 6937 1781 6947
rect 1831 6937 1871 6947
rect 1911 6937 1981 6947
rect 1991 6937 2051 6947
rect 2211 6937 2231 6947
rect 981 6927 1771 6937
rect 741 6917 971 6927
rect 751 6897 971 6917
rect 741 6887 971 6897
rect 731 6852 971 6887
rect 981 6917 1621 6927
rect 1641 6917 1771 6927
rect 1821 6917 1861 6937
rect 1901 6927 2041 6937
rect 2061 6927 2081 6937
rect 1891 6917 2031 6927
rect 2061 6917 2071 6927
rect 2121 6917 2141 6937
rect 2191 6927 2231 6937
rect 2271 6936 2291 6947
rect 2321 6937 2351 6947
rect 2431 6937 2501 6947
rect 2271 6927 2301 6936
rect 2311 6927 2341 6937
rect 2401 6927 2501 6937
rect 2551 6937 2571 6947
rect 2651 6937 2691 6947
rect 2871 6937 2881 6947
rect 2511 6927 2532 6930
rect 2551 6927 2561 6937
rect 2621 6927 2671 6937
rect 2871 6927 2891 6937
rect 2191 6917 2261 6927
rect 2291 6917 2331 6927
rect 2391 6917 2532 6927
rect 2541 6917 2561 6927
rect 2611 6917 2651 6927
rect 2821 6917 2841 6927
rect 2881 6917 2891 6927
rect 981 6897 1601 6917
rect 1631 6907 1781 6917
rect 1801 6907 1811 6917
rect 981 6887 1591 6897
rect 1631 6887 1771 6907
rect 1791 6897 1811 6907
rect 1821 6907 1851 6917
rect 1881 6907 1931 6917
rect 1941 6907 2031 6917
rect 2051 6907 2081 6917
rect 2101 6907 2261 6917
rect 2281 6907 2331 6917
rect 2401 6907 2561 6917
rect 2591 6907 2651 6917
rect 2811 6907 2831 6917
rect 1821 6897 1841 6907
rect 1871 6897 2071 6907
rect 1791 6887 1841 6897
rect 1861 6887 2011 6897
rect 2021 6887 2071 6897
rect 2091 6906 2253 6907
rect 2091 6897 2241 6906
rect 2271 6897 2331 6907
rect 2391 6897 2571 6907
rect 2581 6897 2661 6907
rect 2721 6897 2751 6907
rect 2811 6897 2821 6907
rect 2091 6894 2231 6897
rect 2091 6887 2229 6894
rect 2261 6887 2751 6897
rect 981 6877 1601 6887
rect 1621 6877 1761 6887
rect 1781 6877 1831 6887
rect 981 6867 1591 6877
rect 1621 6867 1731 6877
rect 1741 6867 1761 6877
rect 981 6857 1581 6867
rect 1641 6857 1721 6867
rect 1771 6857 1831 6877
rect 1851 6877 1991 6887
rect 2021 6877 2221 6887
rect 2251 6877 2291 6887
rect 1851 6867 1881 6877
rect 1851 6857 1861 6867
rect 1891 6857 1981 6877
rect 2011 6867 2221 6877
rect 2231 6867 2291 6877
rect 2311 6877 2621 6887
rect 2631 6877 2731 6887
rect 2881 6877 2931 6887
rect 2311 6867 2711 6877
rect 2761 6867 2781 6877
rect 2881 6867 2921 6877
rect 1991 6857 2711 6867
rect 2751 6857 2781 6867
rect 2831 6857 2851 6867
rect 731 6837 781 6852
rect 791 6847 971 6852
rect 991 6847 1571 6857
rect 801 6837 961 6847
rect 991 6837 1561 6847
rect 1641 6837 1711 6857
rect 1761 6847 1831 6857
rect 1891 6847 1931 6857
rect 1971 6847 2781 6857
rect 2811 6847 2851 6857
rect 2931 6847 2961 6857
rect 1761 6837 1821 6847
rect 1891 6837 1921 6847
rect 1961 6837 2841 6847
rect 2921 6837 2961 6847
rect 721 6827 961 6837
rect 981 6827 1551 6837
rect 1651 6827 1701 6837
rect 721 6817 1361 6827
rect 1391 6817 1401 6827
rect 1491 6817 1541 6827
rect 1651 6817 1671 6827
rect 1761 6822 1801 6837
rect 1881 6827 1901 6837
rect 1941 6827 2701 6837
rect 2711 6827 2841 6837
rect 1771 6817 1801 6822
rect 1941 6817 2851 6827
rect 2891 6817 2901 6827
rect 721 6797 781 6817
rect 791 6807 1341 6817
rect 1771 6807 1791 6817
rect 1941 6807 2081 6817
rect 791 6797 1321 6807
rect 1921 6797 1971 6807
rect 1991 6797 2081 6807
rect 2091 6807 2871 6817
rect 2091 6797 2861 6807
rect 751 6787 1261 6797
rect 1281 6787 1311 6797
rect 1921 6787 1961 6797
rect 1991 6787 2121 6797
rect 2131 6787 2171 6797
rect 2191 6787 2781 6797
rect 761 6777 1251 6787
rect 1731 6777 1741 6787
rect 1921 6777 1931 6787
rect 1991 6777 2041 6787
rect 2071 6777 2121 6787
rect 2141 6777 2161 6787
rect 2191 6777 2321 6787
rect 761 6767 1211 6777
rect 1221 6767 1231 6777
rect 1991 6768 2011 6777
rect 1992 6767 2011 6768
rect 2081 6767 2121 6777
rect 2201 6767 2211 6777
rect 2251 6767 2321 6777
rect 2331 6777 2781 6787
rect 2801 6787 2841 6797
rect 2801 6777 2831 6787
rect 2911 6777 2931 6787
rect 2331 6767 2831 6777
rect 761 6757 1181 6767
rect 1992 6757 2001 6767
rect 2081 6757 2091 6767
rect 2101 6757 2111 6767
rect 2251 6757 2844 6767
rect 2881 6757 2891 6767
rect 761 6747 1161 6757
rect 2261 6747 2371 6757
rect 2391 6747 2841 6757
rect 2871 6756 2901 6757
rect 2861 6747 2901 6756
rect 761 6737 1131 6747
rect 2251 6737 2941 6747
rect 761 6727 1111 6737
rect 2251 6727 2971 6737
rect 721 6707 731 6727
rect 761 6717 1101 6727
rect 2241 6717 2981 6727
rect 751 6707 1081 6717
rect 2231 6707 2301 6717
rect 2341 6707 2451 6717
rect 2491 6707 2851 6717
rect 2881 6707 2901 6717
rect 2961 6707 2982 6717
rect 741 6697 1071 6707
rect 2241 6697 2251 6707
rect 2341 6697 2421 6707
rect 2481 6697 2831 6707
rect 2841 6697 2871 6707
rect 2891 6697 2901 6707
rect 741 6687 891 6697
rect 961 6687 1031 6697
rect 2201 6687 2231 6697
rect 2321 6687 2411 6697
rect 2461 6687 2881 6697
rect 731 6677 861 6687
rect 2191 6677 2211 6687
rect 2311 6677 2391 6687
rect 741 6667 851 6677
rect 2291 6667 2371 6677
rect 2421 6667 2441 6677
rect 2451 6667 2891 6687
rect 2931 6677 2941 6687
rect 751 6657 831 6667
rect 2421 6657 2901 6667
rect 761 6647 821 6657
rect 2411 6647 2881 6657
rect 761 6627 811 6647
rect 2401 6637 2861 6647
rect 2311 6627 2341 6637
rect 2361 6627 2411 6637
rect 2471 6627 2871 6637
rect 751 6617 791 6627
rect 2281 6617 2421 6627
rect 2491 6617 2881 6627
rect 761 6607 781 6617
rect 2280 6607 2481 6617
rect 2521 6607 2881 6617
rect 2241 6606 2259 6607
rect 2241 6597 2271 6606
rect 2281 6597 2501 6607
rect 2531 6597 2891 6607
rect 761 6587 771 6597
rect 2251 6587 2261 6597
rect 2311 6587 2911 6597
rect 2331 6577 2911 6587
rect 2321 6557 2331 6567
rect 2351 6557 2861 6577
rect 2883 6567 2931 6577
rect 2271 6547 2441 6557
rect 2461 6547 2861 6557
rect 2871 6552 2907 6567
rect 2951 6557 2971 6577
rect 2871 6547 2901 6552
rect 2281 6537 2531 6547
rect 2541 6537 2901 6547
rect 3001 6537 3021 6567
rect 2251 6527 2261 6537
rect 2291 6527 2831 6537
rect 2841 6527 2901 6537
rect 3031 6527 3051 6537
rect 2291 6517 2821 6527
rect 2841 6517 2911 6527
rect 3031 6517 3061 6527
rect 2301 6507 2911 6517
rect 2311 6497 2841 6507
rect 2221 6487 2231 6497
rect 2251 6487 2361 6497
rect 2281 6477 2361 6487
rect 2391 6477 2791 6497
rect 2811 6487 2851 6497
rect 2861 6487 2911 6507
rect 2841 6477 2921 6487
rect 2291 6467 2381 6477
rect 2391 6467 2801 6477
rect 2851 6467 2871 6477
rect 2911 6467 2941 6477
rect 2311 6447 2811 6467
rect 2961 6456 2982 6468
rect 2971 6447 2981 6456
rect 2321 6437 2821 6447
rect 2891 6437 2911 6447
rect 2971 6437 2991 6447
rect 701 6427 711 6437
rect 2321 6427 2801 6437
rect 2891 6427 2921 6437
rect 2321 6417 2351 6427
rect 2361 6417 2781 6427
rect 2791 6417 2811 6427
rect 2321 6407 2341 6417
rect 2381 6407 2771 6417
rect 2801 6407 2811 6417
rect 2901 6407 2921 6427
rect 2971 6417 3011 6437
rect 2991 6407 3011 6417
rect 2331 6397 2351 6407
rect 2391 6397 2771 6407
rect 2341 6387 2361 6397
rect 2391 6387 2781 6397
rect 2831 6387 2841 6397
rect 2961 6387 2971 6397
rect 2261 6377 2271 6387
rect 2351 6377 2371 6387
rect 2401 6377 2561 6387
rect 2351 6357 2381 6377
rect 2411 6367 2561 6377
rect 2571 6367 2581 6377
rect 2591 6367 2791 6387
rect 2431 6357 2581 6367
rect 2601 6357 2791 6367
rect 2031 6337 2041 6357
rect 2291 6347 2301 6357
rect 2331 6347 2391 6357
rect 2441 6347 2591 6357
rect 2611 6347 2791 6357
rect 2941 6347 2951 6367
rect 2291 6337 2311 6347
rect 2301 6327 2311 6337
rect 2341 6337 2401 6347
rect 2431 6337 2471 6347
rect 2501 6337 2561 6347
rect 2571 6337 2801 6347
rect 2341 6327 2411 6337
rect 2421 6327 2471 6337
rect 2141 6297 2151 6307
rect 2271 6306 2281 6327
rect 2341 6317 2401 6327
rect 2421 6317 2431 6327
rect 2331 6307 2401 6317
rect 2461 6307 2481 6327
rect 2511 6317 2521 6337
rect 2531 6327 2561 6337
rect 2581 6327 2611 6337
rect 2541 6318 2561 6327
rect 2541 6307 2571 6318
rect 2591 6317 2611 6327
rect 2631 6327 2811 6337
rect 2631 6317 2821 6327
rect 2591 6307 2621 6317
rect 2641 6307 2721 6317
rect 2741 6307 2821 6317
rect 2871 6307 2881 6337
rect 2951 6327 2961 6337
rect 2271 6297 2292 6306
rect 2311 6297 2411 6307
rect 2141 6287 2161 6297
rect 2281 6287 2411 6297
rect 2451 6287 2481 6307
rect 2550 6306 2571 6307
rect 2561 6297 2571 6306
rect 2601 6297 2671 6307
rect 2551 6287 2671 6297
rect 2691 6297 2731 6307
rect 2742 6297 2831 6307
rect 2691 6287 2751 6297
rect 2761 6287 2831 6297
rect 2271 6277 2301 6287
rect 2321 6277 2421 6287
rect 2451 6277 2491 6287
rect 2551 6277 2841 6287
rect 2971 6277 2981 6285
rect 2161 6276 2171 6277
rect 2160 6264 2181 6276
rect 2281 6267 2301 6277
rect 2311 6267 2341 6277
rect 2171 6257 2181 6264
rect 2111 6237 2121 6247
rect 2171 6237 2191 6257
rect 2221 6237 2251 6257
rect 2001 6227 2011 6237
rect 2111 6227 2131 6237
rect 2111 6217 2141 6227
rect 2181 6217 2201 6237
rect 2041 6207 2051 6217
rect 2101 6207 2151 6217
rect 2171 6207 2201 6217
rect 2231 6217 2251 6237
rect 2271 6247 2341 6267
rect 2361 6257 2421 6277
rect 2461 6267 2501 6277
rect 2551 6267 2641 6277
rect 2651 6267 2701 6277
rect 2721 6267 2841 6277
rect 2461 6257 2511 6267
rect 2541 6257 2641 6267
rect 2661 6257 2701 6267
rect 2361 6247 2431 6257
rect 2461 6247 2521 6257
rect 2541 6247 2581 6257
rect 2271 6227 2351 6247
rect 2361 6237 2441 6247
rect 2461 6237 2531 6247
rect 2556 6246 2577 6247
rect 2561 6237 2571 6246
rect 2591 6237 2631 6257
rect 2261 6217 2351 6227
rect 2371 6227 2451 6237
rect 2461 6227 2541 6237
rect 2561 6227 2631 6237
rect 2371 6217 2551 6227
rect 2571 6217 2631 6227
rect 2671 6247 2701 6257
rect 2731 6257 2841 6267
rect 2961 6257 3001 6277
rect 2731 6247 2831 6257
rect 2671 6227 2711 6247
rect 2751 6237 2831 6247
rect 2881 6247 2891 6257
rect 2951 6247 3001 6257
rect 2751 6227 2841 6237
rect 2851 6227 2861 6237
rect 2881 6227 2901 6247
rect 2951 6237 2991 6247
rect 2951 6227 2981 6237
rect 2671 6217 2681 6227
rect 2701 6217 2721 6227
rect 2761 6217 2861 6227
rect 2231 6207 2351 6217
rect 2381 6207 2561 6217
rect 2581 6207 2641 6217
rect 2711 6207 2741 6217
rect 2771 6207 2871 6217
rect 1951 6197 1971 6207
rect 2031 6197 2061 6207
rect 2081 6197 2091 6207
rect 2101 6197 2361 6207
rect 2381 6197 2521 6207
rect 2531 6197 2561 6207
rect 2591 6197 2661 6207
rect 2721 6197 2741 6207
rect 2781 6197 2871 6207
rect 2891 6207 2901 6227
rect 2961 6217 2991 6227
rect 2011 6187 2021 6197
rect 2041 6187 2201 6197
rect 2221 6187 2671 6197
rect 2701 6187 2751 6197
rect 2781 6189 2881 6197
rect 2041 6177 2211 6187
rect 2231 6177 2681 6187
rect 2701 6177 2761 6187
rect 2793 6177 2881 6189
rect 2031 6167 2091 6177
rect 2031 6157 2041 6167
rect 2021 6147 2041 6157
rect 2061 6157 2091 6167
rect 2101 6157 2211 6177
rect 2241 6167 2411 6177
rect 2251 6157 2411 6167
rect 2421 6157 2681 6177
rect 2061 6147 2221 6157
rect 2251 6147 2681 6157
rect 2711 6165 2781 6177
rect 2802 6167 2881 6177
rect 2891 6177 2911 6207
rect 2971 6197 2991 6217
rect 2971 6187 3001 6197
rect 2891 6167 2921 6177
rect 2711 6147 2791 6165
rect 2821 6147 2921 6167
rect 2021 6137 2231 6147
rect 2241 6137 2541 6147
rect 2571 6137 2691 6147
rect 2711 6137 2941 6147
rect 1251 6127 1551 6137
rect 2021 6127 2551 6137
rect 2561 6127 2951 6137
rect 1191 6117 1611 6127
rect 2011 6117 2171 6127
rect 2181 6117 2391 6127
rect 1091 6107 1661 6117
rect 2071 6107 2161 6117
rect 2211 6107 2381 6117
rect 1051 6097 1691 6107
rect 2081 6097 2161 6107
rect 2181 6097 2381 6107
rect 2411 6107 2951 6127
rect 2411 6097 2971 6107
rect 781 6087 801 6097
rect 1021 6087 1731 6097
rect 2091 6087 2171 6097
rect 2181 6087 2361 6097
rect 2421 6087 2971 6097
rect 761 6077 851 6087
rect 1011 6077 1571 6087
rect 1641 6077 1771 6087
rect 2091 6077 2191 6087
rect 711 6067 851 6077
rect 991 6067 1571 6077
rect 1661 6067 1811 6077
rect 2071 6067 2191 6077
rect 2221 6077 2361 6087
rect 2431 6077 2951 6087
rect 2221 6067 2391 6077
rect 2421 6067 2941 6077
rect 651 6057 871 6067
rect 991 6057 1581 6067
rect 1651 6057 1881 6067
rect 2081 6057 2621 6067
rect 2641 6057 2701 6067
rect 2721 6057 2941 6067
rect 561 6047 871 6057
rect 501 6037 871 6047
rect 1001 6047 1601 6057
rect 1611 6047 1931 6057
rect 2091 6047 2941 6057
rect 1001 6037 1971 6047
rect 2091 6037 2311 6047
rect 2328 6039 2501 6047
rect 2328 6037 2481 6039
rect 2511 6037 2651 6047
rect 2661 6037 2941 6047
rect 461 6027 861 6037
rect 441 6017 861 6027
rect 1001 6027 2051 6037
rect 2081 6027 2352 6037
rect 1001 6017 2251 6027
rect 2291 6017 2361 6027
rect 2381 6017 2481 6037
rect 2541 6027 2931 6037
rect 2491 6017 2511 6027
rect 2551 6017 2931 6027
rect 421 6007 861 6017
rect 911 6007 921 6017
rect 961 6007 971 6017
rect 991 6007 1691 6017
rect 1791 6007 2261 6017
rect 2291 6007 2301 6017
rect 2311 6007 2431 6017
rect 2451 6007 2531 6017
rect 2571 6007 2771 6017
rect 2781 6007 2931 6017
rect 401 5997 871 6007
rect 911 5997 1671 6007
rect 1861 5997 2271 6007
rect 2281 5997 2301 6007
rect 2321 5997 2441 6007
rect 2461 5997 2531 6007
rect 2581 5997 2951 6007
rect 371 5987 1651 5997
rect 1951 5987 2361 5997
rect 2391 5987 2541 5997
rect 351 5977 941 5987
rect 951 5977 1641 5987
rect 2021 5977 2551 5987
rect 2591 5977 2931 5997
rect 2941 5987 2951 5997
rect 341 5967 901 5977
rect 961 5967 1631 5977
rect 2081 5967 2561 5977
rect 321 5957 891 5967
rect 311 5947 891 5957
rect 291 5937 891 5947
rect 291 5927 311 5937
rect 341 5927 891 5937
rect 291 5917 301 5927
rect 341 5907 821 5927
rect 331 5897 821 5907
rect 831 5897 891 5927
rect 981 5957 1041 5967
rect 1051 5957 1631 5967
rect 2131 5957 2561 5967
rect 2601 5967 2931 5977
rect 2941 5967 2951 5977
rect 2601 5957 2951 5967
rect 981 5947 1621 5957
rect 2181 5947 2941 5957
rect 981 5937 1591 5947
rect 2201 5946 2931 5947
rect 2201 5937 2461 5946
rect 2481 5937 2931 5946
rect 981 5897 1041 5937
rect 1051 5897 1581 5937
rect 2211 5927 2471 5937
rect 2491 5927 2931 5937
rect 2211 5917 2321 5927
rect 2331 5917 2481 5927
rect 2501 5917 2551 5927
rect 2561 5917 2921 5927
rect 2211 5907 2491 5917
rect 2511 5907 2921 5917
rect 2171 5897 2181 5907
rect 2211 5897 2501 5907
rect 2521 5897 2921 5907
rect 311 5887 881 5897
rect 291 5867 881 5887
rect 991 5867 1041 5897
rect 291 5857 871 5867
rect 321 5847 871 5857
rect 1001 5847 1041 5867
rect 1061 5887 1581 5897
rect 2111 5887 2511 5897
rect 2521 5887 2571 5897
rect 2661 5887 2921 5897
rect 331 5837 861 5847
rect 341 5827 861 5837
rect 1001 5827 1051 5847
rect 341 5817 421 5827
rect 431 5817 831 5827
rect 841 5817 851 5827
rect 341 5807 831 5817
rect 371 5797 831 5807
rect 1011 5807 1051 5827
rect 1061 5817 1591 5887
rect 2061 5877 2541 5887
rect 2681 5877 2911 5887
rect 2051 5857 2521 5877
rect 2701 5867 2911 5877
rect 2711 5857 2911 5867
rect 2051 5847 2511 5857
rect 2721 5847 2901 5857
rect 2061 5837 2151 5847
rect 2191 5837 2491 5847
rect 2731 5837 2901 5847
rect 2081 5827 2091 5837
rect 2211 5827 2351 5837
rect 2371 5827 2451 5837
rect 2741 5827 2901 5837
rect 2221 5817 2331 5827
rect 2371 5817 2401 5827
rect 2421 5817 2451 5827
rect 1011 5797 1061 5807
rect 391 5767 821 5797
rect 1021 5787 1061 5797
rect 1071 5787 1591 5817
rect 1021 5777 1051 5787
rect 1081 5777 1591 5787
rect 2251 5797 2321 5817
rect 2381 5807 2391 5817
rect 2751 5807 2901 5827
rect 2641 5797 2651 5807
rect 2761 5797 2901 5807
rect 401 5757 411 5767
rect 421 5757 821 5767
rect 1081 5757 1581 5777
rect 2251 5767 2281 5797
rect 2291 5787 2321 5797
rect 2671 5787 2681 5797
rect 2771 5787 2901 5797
rect 2291 5777 2311 5787
rect 2531 5777 2561 5787
rect 2671 5777 2701 5787
rect 2781 5777 2901 5787
rect 2231 5757 2281 5767
rect 2521 5757 2551 5777
rect 2681 5767 2711 5777
rect 2781 5767 2891 5777
rect 2691 5757 2721 5767
rect 2791 5757 2891 5767
rect 401 5737 831 5757
rect 401 5697 821 5737
rect 1061 5727 1071 5736
rect 1061 5717 1081 5727
rect 1091 5717 1581 5757
rect 1621 5747 1641 5757
rect 2231 5747 2251 5757
rect 2141 5737 2161 5747
rect 2121 5727 2161 5737
rect 2221 5737 2251 5747
rect 2221 5727 2231 5737
rect 2511 5727 2551 5757
rect 2701 5747 2731 5757
rect 2681 5737 2741 5747
rect 2791 5737 2881 5757
rect 2721 5727 2741 5737
rect 2121 5717 2151 5727
rect 2211 5717 2231 5727
rect 2701 5717 2741 5727
rect 2801 5727 2831 5737
rect 2841 5727 2881 5737
rect 1071 5707 1081 5717
rect 1101 5697 1581 5717
rect 2131 5707 2151 5717
rect 2181 5707 2201 5717
rect 2171 5697 2201 5707
rect 2711 5707 2751 5717
rect 2801 5707 2821 5727
rect 2861 5717 2871 5727
rect 401 5677 811 5697
rect 1111 5677 1571 5697
rect 2171 5687 2191 5697
rect 401 5647 801 5677
rect 1121 5667 1561 5677
rect 1131 5657 1561 5667
rect 2481 5667 2501 5677
rect 2711 5667 2741 5707
rect 2481 5657 2521 5667
rect 1131 5647 1551 5657
rect 411 5617 791 5647
rect 1141 5637 1551 5647
rect 2471 5647 2541 5657
rect 2721 5647 2741 5667
rect 2801 5697 2831 5707
rect 2801 5687 2861 5697
rect 2801 5677 2831 5687
rect 2841 5677 2851 5687
rect 2801 5647 2851 5677
rect 2471 5637 2551 5647
rect 2721 5637 2751 5647
rect 1151 5617 1541 5637
rect 2471 5627 2571 5637
rect 2481 5617 2571 5627
rect 2721 5617 2741 5637
rect 2801 5627 2841 5647
rect 421 5607 791 5617
rect 1171 5607 1531 5617
rect 2481 5607 2581 5617
rect 421 5587 781 5607
rect 1181 5597 1521 5607
rect 1191 5587 1511 5597
rect 431 5567 771 5587
rect 1091 5577 1121 5587
rect 1211 5577 1491 5587
rect 2481 5577 2521 5607
rect 2541 5597 2561 5607
rect 2721 5597 2731 5617
rect 2801 5597 2811 5627
rect 2821 5617 2841 5627
rect 2541 5577 2551 5597
rect 2791 5587 2811 5597
rect 1041 5567 1051 5577
rect 1081 5567 1131 5577
rect 1231 5567 1471 5577
rect 2491 5567 2511 5577
rect 2791 5567 2821 5587
rect 441 5557 771 5567
rect 1081 5557 1141 5567
rect 1231 5557 1451 5567
rect 2781 5557 2801 5567
rect 451 5537 761 5557
rect 1081 5547 1161 5557
rect 1211 5547 1401 5557
rect 2781 5547 2791 5557
rect 2811 5547 2821 5567
rect 1091 5537 1171 5547
rect 1201 5537 1261 5547
rect 2771 5537 2791 5547
rect 461 5527 751 5537
rect 471 5517 741 5527
rect 1101 5517 1251 5537
rect 2431 5517 2441 5527
rect 481 5507 731 5517
rect 1101 5507 1211 5517
rect 1221 5507 1251 5517
rect 2451 5507 2471 5517
rect 2761 5507 2791 5537
rect 491 5497 731 5507
rect 1111 5497 1211 5507
rect 2461 5497 2471 5507
rect 2601 5497 2621 5507
rect 2751 5497 2781 5507
rect 511 5487 721 5497
rect 1121 5487 1231 5497
rect 551 5477 631 5487
rect 691 5477 721 5487
rect 1131 5477 1231 5487
rect 2741 5477 2781 5497
rect 701 5467 711 5477
rect 1121 5467 1241 5477
rect 1131 5457 1251 5467
rect 2731 5457 2771 5477
rect 1131 5447 1261 5457
rect 761 5437 781 5447
rect 1131 5437 1271 5447
rect 2721 5437 2771 5457
rect 761 5427 791 5437
rect 1121 5427 1281 5437
rect 2711 5427 2761 5437
rect 771 5417 811 5427
rect 1121 5417 1291 5427
rect 771 5407 821 5417
rect 941 5407 1051 5417
rect 1111 5407 1291 5417
rect 2701 5407 2761 5427
rect 781 5397 831 5407
rect 901 5397 1071 5407
rect 1101 5397 1311 5407
rect 2691 5397 2751 5407
rect 781 5387 851 5397
rect 871 5387 1311 5397
rect 2681 5387 2751 5397
rect 781 5377 861 5387
rect 871 5377 1321 5387
rect 2671 5377 2751 5387
rect 781 5367 1321 5377
rect 2661 5367 2741 5377
rect 751 5357 1131 5367
rect 1161 5357 1321 5367
rect 2651 5357 2741 5367
rect 751 5347 1111 5357
rect 1161 5347 1331 5357
rect 2641 5347 2731 5357
rect 741 5337 891 5347
rect 901 5337 1111 5347
rect 1181 5337 1331 5347
rect 2371 5337 2411 5347
rect 2631 5337 2731 5347
rect 741 5327 1131 5337
rect 1211 5328 1331 5337
rect 1233 5327 1331 5328
rect 2621 5327 2721 5337
rect 741 5307 841 5327
rect 851 5317 1131 5327
rect 1241 5317 1331 5327
rect 2611 5317 2721 5327
rect 611 5287 631 5307
rect 741 5297 831 5307
rect 871 5297 1051 5317
rect 1071 5307 1131 5317
rect 1233 5316 1331 5317
rect 1221 5307 1331 5316
rect 1361 5307 1371 5317
rect 2611 5307 2711 5317
rect 1061 5297 1121 5307
rect 1251 5297 1341 5307
rect 741 5287 811 5297
rect 731 5277 811 5287
rect 871 5287 1111 5297
rect 1261 5287 1351 5297
rect 2301 5287 2331 5297
rect 871 5277 1101 5287
rect 1271 5277 1361 5287
rect 2291 5277 2331 5287
rect 2601 5277 2701 5307
rect 731 5267 801 5277
rect 601 5247 651 5267
rect 611 5237 651 5247
rect 721 5257 791 5267
rect 891 5257 1101 5277
rect 1281 5267 1371 5277
rect 1161 5257 1181 5267
rect 1311 5257 1361 5267
rect 2291 5257 2321 5277
rect 2591 5257 2691 5277
rect 721 5247 781 5257
rect 871 5247 1001 5257
rect 1041 5247 1051 5257
rect 1061 5247 1101 5257
rect 2291 5247 2311 5257
rect 2591 5247 2681 5257
rect 721 5237 771 5247
rect 601 5227 651 5237
rect 731 5227 771 5237
rect 871 5237 991 5247
rect 1071 5237 1101 5247
rect 2581 5237 2681 5247
rect 871 5227 1001 5237
rect 1091 5227 1111 5237
rect 2581 5227 2671 5237
rect 601 5217 661 5227
rect 591 5207 661 5217
rect 721 5217 761 5227
rect 721 5207 751 5217
rect 871 5207 981 5227
rect 561 5187 571 5207
rect 581 5187 671 5207
rect 721 5197 741 5207
rect 861 5197 981 5207
rect 2571 5207 2661 5227
rect 2571 5197 2631 5207
rect 2641 5197 2651 5207
rect 591 5157 671 5187
rect 861 5187 971 5197
rect 861 5177 951 5187
rect 2561 5177 2631 5197
rect 901 5167 931 5177
rect 601 5147 671 5157
rect 2551 5157 2631 5177
rect 2551 5147 2621 5157
rect 601 5117 681 5147
rect 971 5137 1041 5147
rect 2551 5137 2611 5147
rect 841 5127 871 5137
rect 951 5127 1081 5137
rect 841 5117 911 5127
rect 931 5117 1121 5127
rect 2541 5117 2611 5137
rect 611 5097 681 5117
rect 831 5107 1151 5117
rect 821 5097 1181 5107
rect 2541 5097 2591 5117
rect 621 5087 681 5097
rect 822 5087 1211 5097
rect 641 5077 671 5087
rect 822 5077 1221 5087
rect 1241 5077 1311 5087
rect 2531 5077 2581 5097
rect 822 5076 1351 5077
rect 801 5067 811 5073
rect 821 5067 1351 5076
rect 801 5057 1371 5067
rect 2531 5057 2571 5077
rect 741 5047 751 5057
rect 791 5047 1381 5057
rect 731 5037 761 5047
rect 791 5037 1391 5047
rect 2521 5037 2561 5057
rect 731 5027 1051 5037
rect 1121 5027 1141 5037
rect 1151 5027 1411 5037
rect 731 5017 1001 5027
rect 1191 5017 1211 5027
rect 1241 5017 1411 5027
rect 731 5007 961 5017
rect 1271 5007 1421 5017
rect 2521 5007 2551 5037
rect 731 4997 843 5007
rect 873 4997 951 5007
rect 1331 4997 1431 5007
rect 731 4987 841 4997
rect 891 4987 921 4997
rect 1351 4987 1411 4997
rect 1421 4987 1431 4997
rect 731 4967 831 4987
rect 891 4977 901 4987
rect 881 4967 901 4977
rect 1371 4977 1401 4987
rect 1421 4977 1441 4987
rect 2511 4977 2541 5007
rect 1371 4967 1451 4977
rect 2511 4967 2531 4977
rect 731 4957 821 4967
rect 741 4947 801 4957
rect 881 4947 891 4967
rect 1021 4957 1031 4967
rect 1391 4957 1451 4967
rect 911 4947 951 4957
rect 1401 4947 1451 4957
rect 741 4937 781 4947
rect 881 4937 971 4947
rect 1411 4937 1451 4947
rect 751 4907 781 4937
rect 851 4927 981 4937
rect 1431 4927 1451 4937
rect 2501 4957 2531 4967
rect 2501 4937 2521 4957
rect 841 4917 981 4927
rect 2501 4917 2511 4937
rect 851 4907 981 4917
rect 761 4897 771 4907
rect 861 4897 1001 4907
rect 851 4887 1031 4897
rect 2491 4887 2501 4907
rect 851 4867 1051 4887
rect 841 4857 1061 4867
rect 1091 4857 1121 4867
rect 851 4847 1171 4857
rect 611 4837 631 4847
rect 651 4837 661 4847
rect 851 4837 1191 4847
rect 861 4817 1221 4837
rect 521 4797 591 4817
rect 851 4807 1231 4817
rect 851 4797 1241 4807
rect 531 4787 571 4797
rect 851 4787 1251 4797
rect 531 4777 601 4787
rect 731 4777 741 4787
rect 851 4777 1261 4787
rect 541 4757 611 4777
rect 861 4767 1261 4777
rect 861 4757 1251 4767
rect 571 4747 601 4757
rect 851 4747 1231 4757
rect 321 4737 331 4747
rect 551 4737 601 4747
rect 861 4737 1221 4747
rect 301 4727 331 4737
rect 531 4697 591 4737
rect 861 4728 1081 4737
rect 861 4727 1065 4728
rect 1121 4727 1221 4737
rect 871 4719 1065 4727
rect 871 4717 1041 4719
rect 1141 4717 1191 4727
rect 881 4707 1041 4717
rect 891 4697 931 4707
rect 971 4697 1041 4707
rect 531 4677 571 4697
rect 891 4687 911 4697
rect 981 4687 1031 4697
rect 1051 4687 1061 4707
rect 531 4667 591 4677
rect 531 4657 601 4667
rect 971 4657 1041 4687
rect 461 4647 511 4657
rect 521 4647 611 4657
rect 801 4647 831 4657
rect 451 4637 611 4647
rect 811 4637 831 4647
rect 441 4627 611 4637
rect 821 4627 841 4637
rect 971 4627 1051 4657
rect 441 4617 511 4627
rect 531 4617 641 4627
rect 731 4617 771 4627
rect 971 4617 1061 4627
rect 441 4597 491 4617
rect 541 4608 651 4617
rect 541 4607 630 4608
rect 961 4607 1071 4617
rect 551 4597 630 4607
rect 951 4597 1081 4607
rect 561 4577 611 4597
rect 791 4587 821 4597
rect 801 4577 821 4587
rect 561 4567 571 4577
rect 581 4567 601 4577
rect 591 4547 601 4567
rect 831 4557 841 4577
rect 971 4567 1091 4597
rect 921 4557 1111 4567
rect 931 4547 1121 4557
rect 921 4537 1121 4547
rect 921 4527 1201 4537
rect 921 4517 1211 4527
rect 1231 4517 1241 4527
rect 841 4507 861 4517
rect 921 4507 1271 4517
rect 781 4506 792 4507
rect 781 4497 811 4506
rect 801 4487 811 4497
rect 921 4497 1281 4507
rect 921 4487 1311 4497
rect 921 4477 1341 4487
rect 921 4467 1351 4477
rect 931 4447 1371 4467
rect 1401 4457 1431 4467
rect 1411 4447 1431 4457
rect 901 4437 921 4447
rect 941 4437 1381 4447
rect 1761 4437 1771 4447
rect 931 4427 1391 4437
rect 1421 4427 1431 4437
rect 1571 4427 1601 4437
rect 1611 4427 1671 4437
rect 1731 4427 1751 4437
rect 2481 4427 2491 4437
rect 861 4417 871 4427
rect 931 4417 1371 4427
rect 1401 4417 1471 4427
rect 1531 4417 1771 4427
rect 801 4397 811 4417
rect 861 4407 881 4417
rect 971 4407 1361 4417
rect 1001 4397 1361 4407
rect 1391 4407 1491 4417
rect 1511 4407 1771 4417
rect 2471 4407 2501 4427
rect 1391 4397 1741 4407
rect 2471 4397 2481 4407
rect 791 4387 811 4397
rect 831 4387 851 4397
rect 871 4387 891 4397
rect 1011 4387 1741 4397
rect 781 4377 921 4387
rect 1001 4377 1751 4387
rect 2461 4377 2481 4397
rect 2511 4387 2531 4397
rect 2521 4377 2531 4387
rect 771 4367 941 4377
rect 771 4357 851 4367
rect 881 4357 941 4367
rect 991 4357 1201 4377
rect 1221 4367 1281 4377
rect 1291 4367 1751 4377
rect 2471 4367 2491 4377
rect 751 4347 801 4357
rect 831 4347 951 4357
rect 981 4347 1201 4357
rect 1231 4347 1301 4367
rect 1321 4357 1771 4367
rect 2471 4357 2511 4367
rect 1331 4347 1791 4357
rect 411 4337 421 4347
rect 711 4337 811 4347
rect 491 4317 501 4337
rect 621 4327 811 4337
rect 611 4317 811 4327
rect 821 4337 941 4347
rect 971 4337 1201 4347
rect 1251 4337 1301 4347
rect 821 4327 1221 4337
rect 1261 4327 1311 4337
rect 1341 4327 1801 4347
rect 2481 4337 2511 4357
rect 2491 4327 2511 4337
rect 821 4317 1231 4327
rect 441 4307 501 4317
rect 601 4307 721 4317
rect 431 4297 501 4307
rect 591 4297 721 4307
rect 731 4307 1181 4317
rect 731 4297 751 4307
rect 781 4297 1171 4307
rect 1191 4297 1231 4317
rect 1261 4317 1321 4327
rect 1331 4317 1811 4327
rect 2501 4317 2511 4327
rect 1261 4307 1351 4317
rect 1381 4307 1811 4317
rect 2471 4307 2481 4317
rect 1271 4297 1351 4307
rect 391 4287 402 4297
rect 441 4287 511 4297
rect 591 4287 741 4297
rect 781 4287 1181 4297
rect 1191 4287 1241 4297
rect 1291 4287 1351 4297
rect 1391 4287 1811 4307
rect 411 4277 521 4287
rect 581 4277 1261 4287
rect 391 4267 531 4277
rect 581 4267 891 4277
rect 901 4267 1201 4277
rect 1211 4267 1261 4277
rect 1301 4277 1361 4287
rect 1391 4277 1801 4287
rect 1301 4267 1371 4277
rect 1381 4267 1811 4277
rect 391 4257 571 4267
rect 581 4257 1201 4267
rect 391 4247 1201 4257
rect 391 4237 811 4247
rect 821 4237 1201 4247
rect 391 4227 841 4237
rect 851 4227 1201 4237
rect 1221 4247 1271 4267
rect 1301 4247 1411 4267
rect 1441 4257 1801 4267
rect 2461 4257 2481 4307
rect 2511 4287 2521 4297
rect 1221 4227 1311 4247
rect 1341 4237 1411 4247
rect 391 4217 831 4227
rect 851 4217 1231 4227
rect 1251 4217 1311 4227
rect 421 4207 821 4217
rect 431 4197 621 4207
rect 631 4197 801 4207
rect 451 4177 581 4197
rect 671 4187 771 4197
rect 841 4187 1231 4217
rect 1261 4207 1311 4217
rect 1351 4227 1411 4237
rect 1451 4247 1791 4257
rect 1451 4237 1781 4247
rect 2461 4237 2491 4257
rect 1451 4227 1791 4237
rect 2461 4227 2501 4237
rect 1351 4217 1811 4227
rect 1261 4197 1321 4207
rect 1351 4197 1471 4217
rect 1511 4197 1811 4217
rect 1261 4187 1371 4197
rect 1401 4187 1471 4197
rect 1521 4187 1831 4197
rect 2461 4187 2511 4227
rect 681 4177 731 4187
rect 741 4177 781 4187
rect 831 4177 1241 4187
rect 1271 4179 1371 4187
rect 1290 4177 1371 4179
rect 461 4167 571 4177
rect 691 4167 731 4177
rect 761 4167 781 4177
rect 821 4167 1251 4177
rect 1301 4167 1371 4177
rect 1411 4177 1481 4187
rect 1511 4177 1831 4187
rect 1411 4167 1491 4177
rect 1511 4167 1541 4177
rect 1561 4167 1831 4177
rect 2451 4177 2501 4187
rect 2451 4167 2491 4177
rect 471 4157 561 4167
rect 761 4157 771 4167
rect 821 4157 1271 4167
rect 541 4147 561 4157
rect 691 4147 701 4157
rect 811 4147 1271 4157
rect 1311 4157 1371 4167
rect 1421 4157 1541 4167
rect 1581 4157 1831 4167
rect 1311 4147 1381 4157
rect 1411 4147 1531 4157
rect 1581 4147 1671 4157
rect 1681 4147 1831 4157
rect 2441 4147 2481 4167
rect 691 4127 721 4147
rect 731 4127 741 4147
rect 811 4137 1281 4147
rect 791 4127 1281 4137
rect 1321 4128 1431 4147
rect 1461 4137 1541 4147
rect 1341 4127 1431 4128
rect 1471 4127 1541 4137
rect 1591 4137 1841 4147
rect 2431 4137 2471 4147
rect 1591 4127 1851 4137
rect 2431 4127 2461 4137
rect 691 4117 701 4127
rect 791 4117 1301 4127
rect 781 4116 1314 4117
rect 781 4107 1321 4116
rect 1361 4107 1431 4127
rect 1481 4117 1551 4127
rect 1581 4117 1621 4127
rect 1631 4117 1861 4127
rect 2421 4117 2451 4127
rect 1481 4107 1611 4117
rect 771 4097 1321 4107
rect 1371 4097 1441 4107
rect 1471 4097 1601 4107
rect 1651 4097 1731 4117
rect 1771 4107 1860 4117
rect 2411 4107 2441 4117
rect 2701 4107 2711 4117
rect 1771 4097 1831 4107
rect 1851 4097 1861 4107
rect 2411 4097 2431 4107
rect 761 4087 1331 4097
rect 701 4077 711 4087
rect 751 4077 1331 4087
rect 1381 4087 1451 4097
rect 1461 4087 1491 4097
rect 1531 4087 1601 4097
rect 1661 4087 1741 4097
rect 1771 4087 1861 4097
rect 2401 4087 2421 4097
rect 1381 4077 1491 4087
rect 611 4067 631 4077
rect 691 4067 711 4077
rect 741 4067 1341 4077
rect 1371 4067 1391 4077
rect 1411 4067 1491 4077
rect 1541 4077 1611 4087
rect 1661 4077 1821 4087
rect 1831 4077 1871 4087
rect 2401 4077 2411 4087
rect 1541 4067 1621 4077
rect 1651 4067 1801 4077
rect 1851 4067 1891 4077
rect 731 4057 1381 4067
rect 591 4047 611 4057
rect 651 4047 1381 4057
rect 1431 4057 1491 4067
rect 1551 4057 1671 4067
rect 1721 4057 1801 4067
rect 1871 4057 1911 4067
rect 1431 4047 1501 4057
rect 1531 4047 1671 4057
rect 571 4037 1301 4047
rect 1321 4037 1391 4047
rect 531 4027 1301 4037
rect 501 4017 1301 4027
rect 1331 4027 1391 4037
rect 1441 4037 1561 4047
rect 1591 4037 1671 4047
rect 1441 4027 1551 4037
rect 1331 4017 1411 4027
rect 1441 4026 1451 4027
rect 1481 4017 1551 4027
rect 1611 4027 1671 4037
rect 1731 4037 1801 4057
rect 1881 4047 1911 4057
rect 1731 4027 1800 4037
rect 1611 4017 1681 4027
rect 1776 4026 1801 4027
rect 1791 4017 1801 4026
rect 461 4007 1311 4017
rect 1341 4007 1441 4017
rect 391 3997 1441 4007
rect 1491 4007 1561 4017
rect 1621 4007 1711 4017
rect 1811 4007 1851 4017
rect 1491 3997 1571 4007
rect 1621 3997 1721 4007
rect 341 3987 1351 3997
rect 1381 3987 1451 3997
rect 311 3977 1351 3987
rect 281 3967 1351 3977
rect 251 3957 1351 3967
rect 1391 3977 1451 3987
rect 1501 3987 1581 3997
rect 1601 3987 1611 3997
rect 1661 3987 1731 3997
rect 1811 3987 1861 4007
rect 1961 3997 1971 4027
rect 2581 4017 2601 4037
rect 2581 4007 2611 4017
rect 2581 3987 2621 4007
rect 1501 3977 1621 3987
rect 1671 3977 1741 3987
rect 1821 3977 1871 3987
rect 1391 3967 1471 3977
rect 1491 3967 1511 3977
rect 1541 3967 1621 3977
rect 1391 3957 1511 3967
rect 221 3947 1371 3957
rect 1381 3947 1511 3957
rect 201 3937 1411 3947
rect 1441 3937 1511 3947
rect 171 3927 1401 3937
rect 1451 3927 1511 3937
rect 1561 3957 1621 3967
rect 1691 3967 1741 3977
rect 1841 3967 1851 3977
rect 2591 3967 2621 3987
rect 1691 3957 1751 3967
rect 1891 3957 1921 3967
rect 2581 3957 2621 3967
rect 1561 3937 1631 3957
rect 1711 3947 1761 3957
rect 1881 3947 1931 3957
rect 1741 3937 1801 3947
rect 1561 3927 1671 3937
rect 1751 3927 1811 3937
rect 1891 3927 1931 3947
rect 2031 3947 2041 3957
rect 2581 3947 2631 3957
rect 2031 3937 2051 3947
rect 2581 3927 2651 3947
rect 121 3917 1411 3927
rect 1451 3917 1531 3927
rect 1611 3917 1681 3927
rect 91 3907 1411 3917
rect 1461 3907 1561 3917
rect 1621 3907 1681 3917
rect 1761 3907 1811 3927
rect 2581 3917 2661 3927
rect 3421 3917 3429 3927
rect 2581 3907 2671 3917
rect 3228 3909 3251 3917
rect 3211 3907 3251 3909
rect 71 3897 1421 3907
rect 1451 3897 1571 3907
rect 45 3877 1471 3897
rect 1511 3887 1571 3897
rect 1631 3897 1691 3907
rect 1771 3897 1811 3907
rect 1631 3887 1701 3897
rect 1821 3887 1861 3897
rect 1511 3877 1581 3887
rect 1641 3877 1731 3887
rect 45 3867 1461 3877
rect 1521 3867 1591 3877
rect 1671 3867 1741 3877
rect 1821 3867 1881 3887
rect 1961 3877 2001 3907
rect 2101 3897 2111 3907
rect 2241 3897 2261 3907
rect 2101 3887 2121 3897
rect 2241 3887 2291 3897
rect 2231 3877 2301 3887
rect 1971 3867 1991 3877
rect 2121 3867 2141 3877
rect 2201 3867 2311 3877
rect 2581 3867 2681 3907
rect 3201 3897 3261 3907
rect 3191 3887 3261 3897
rect 3191 3867 3271 3887
rect 3401 3867 3429 3917
rect 45 3837 1381 3867
rect 1401 3857 1471 3867
rect 1521 3857 1621 3867
rect 1691 3857 1751 3867
rect 1831 3857 1871 3867
rect 2121 3857 2151 3867
rect 2181 3857 2321 3867
rect 2581 3857 2691 3867
rect 2731 3857 2761 3867
rect 3191 3857 3281 3867
rect 1411 3847 1481 3857
rect 1511 3847 1631 3857
rect 1411 3837 1531 3847
rect 1571 3837 1641 3847
rect 1701 3837 1761 3857
rect 1851 3847 1871 3857
rect 2111 3847 2151 3857
rect 2171 3847 2331 3857
rect 2581 3847 2781 3857
rect 3181 3847 3291 3857
rect 3411 3847 3429 3867
rect 1901 3837 1921 3847
rect 2041 3837 2071 3847
rect 2111 3837 2141 3847
rect 2171 3837 2341 3847
rect 2581 3837 2811 3847
rect 3191 3837 3291 3847
rect 45 3827 1391 3837
rect 1411 3827 1521 3837
rect 45 3787 1431 3827
rect 1451 3817 1531 3827
rect 1581 3817 1651 3837
rect 1711 3827 1761 3837
rect 1771 3827 1781 3837
rect 1901 3827 1941 3837
rect 2031 3827 2071 3837
rect 2181 3827 2351 3837
rect 1751 3817 1811 3827
rect 1461 3807 1531 3817
rect 1591 3807 1671 3817
rect 1761 3807 1821 3817
rect 1901 3807 1951 3827
rect 2041 3817 2071 3827
rect 2201 3817 2351 3827
rect 2581 3827 2821 3837
rect 3191 3827 3281 3837
rect 3391 3827 3429 3847
rect 2581 3817 2861 3827
rect 3181 3817 3271 3827
rect 3411 3817 3429 3827
rect 2201 3807 2361 3817
rect 2581 3807 2871 3817
rect 3191 3807 3271 3817
rect 1471 3797 1541 3807
rect 1601 3797 1701 3807
rect 1471 3787 1561 3797
rect 1641 3787 1711 3797
rect 1771 3787 1831 3807
rect 1911 3797 1941 3807
rect 2091 3797 2101 3807
rect 2211 3797 2371 3807
rect 2071 3787 2111 3797
rect 2221 3787 2371 3797
rect 2581 3797 2921 3807
rect 3201 3797 3271 3807
rect 3421 3797 3429 3817
rect 45 3777 1441 3787
rect 1471 3777 1591 3787
rect 45 3767 1451 3777
rect 1471 3767 1491 3777
rect 1521 3767 1591 3777
rect 1651 3777 1711 3787
rect 1781 3777 1831 3787
rect 2001 3777 2011 3787
rect 1651 3767 1721 3777
rect 1811 3767 1841 3777
rect 1851 3767 1871 3777
rect 1991 3767 2021 3777
rect 45 3747 1481 3767
rect 1531 3757 1601 3767
rect 1661 3757 1731 3767
rect 1831 3757 1881 3767
rect 1981 3757 2021 3767
rect 2071 3767 2101 3787
rect 2221 3777 2381 3787
rect 2171 3767 2251 3777
rect 2071 3757 2111 3767
rect 2121 3757 2241 3767
rect 2271 3757 2391 3777
rect 2581 3767 2761 3797
rect 2781 3787 2931 3797
rect 3191 3787 3261 3797
rect 2791 3777 2971 3787
rect 3191 3777 3251 3787
rect 3391 3777 3429 3787
rect 2791 3767 2981 3777
rect 2581 3757 2771 3767
rect 2811 3757 2981 3767
rect 3191 3757 3241 3777
rect 1541 3747 1601 3757
rect 1671 3747 1761 3757
rect 1841 3747 1891 3757
rect 1981 3747 2011 3757
rect 2081 3747 2201 3757
rect 2211 3747 2241 3757
rect 2291 3747 2322 3757
rect 45 3737 1491 3747
rect 1541 3737 1611 3747
rect 1701 3737 1771 3747
rect 1841 3737 1901 3747
rect 2071 3738 2241 3747
rect 2071 3737 2253 3738
rect 45 3727 1501 3737
rect 1551 3727 1651 3737
rect 1711 3727 1781 3737
rect 1851 3727 1891 3737
rect 2031 3727 2171 3737
rect 2181 3727 2201 3737
rect 2231 3729 2253 3737
rect 2301 3735 2322 3747
rect 2331 3747 2401 3757
rect 2581 3747 2781 3757
rect 2331 3737 2341 3747
rect 2231 3727 2262 3729
rect 2311 3727 2321 3735
rect 2351 3727 2411 3747
rect 2581 3737 2791 3747
rect 2581 3727 2811 3737
rect 2821 3727 3011 3757
rect 3191 3747 3251 3757
rect 3051 3727 3071 3747
rect 45 3717 1511 3727
rect 1581 3717 1661 3727
rect 1721 3717 1791 3727
rect 1871 3717 1891 3727
rect 2021 3717 2191 3727
rect 2238 3717 2281 3727
rect 2341 3717 2361 3727
rect 45 3707 1541 3717
rect 1601 3707 1661 3717
rect 1731 3707 1791 3717
rect 45 3697 1551 3707
rect 45 3657 1461 3697
rect 1471 3687 1551 3697
rect 1611 3697 1671 3707
rect 1731 3697 1831 3707
rect 1911 3697 1951 3717
rect 2021 3707 2181 3717
rect 2201 3707 2211 3717
rect 2021 3697 2211 3707
rect 2238 3707 2291 3717
rect 2331 3708 2351 3717
rect 2371 3708 2421 3727
rect 2581 3717 3011 3727
rect 3061 3717 3081 3727
rect 3191 3717 3261 3747
rect 2331 3707 2421 3708
rect 2571 3707 3051 3717
rect 2238 3697 2301 3707
rect 2341 3697 2431 3707
rect 1611 3687 1681 3697
rect 1771 3687 1841 3697
rect 1911 3687 1961 3697
rect 1491 3677 1561 3687
rect 1611 3677 1711 3687
rect 1781 3677 1841 3687
rect 1921 3677 1961 3687
rect 2011 3677 2331 3697
rect 2343 3696 2431 3697
rect 2351 3687 2431 3696
rect 2341 3677 2441 3687
rect 1491 3667 1571 3677
rect 1611 3667 1621 3677
rect 1641 3667 1721 3677
rect 1791 3667 1851 3677
rect 1941 3667 1951 3677
rect 2001 3667 2441 3677
rect 2581 3677 3081 3707
rect 3211 3697 3261 3717
rect 3371 3697 3381 3717
rect 3121 3687 3131 3697
rect 3211 3687 3241 3697
rect 3121 3677 3141 3687
rect 3211 3677 3221 3687
rect 3271 3677 3291 3697
rect 2581 3667 3091 3677
rect 3121 3667 3151 3677
rect 1491 3657 1621 3667
rect 1661 3657 1731 3667
rect 1791 3657 1861 3667
rect 1991 3657 2451 3667
rect 2581 3657 2891 3667
rect 2901 3657 3141 3667
rect 45 3647 1611 3657
rect 1671 3647 1731 3657
rect 1801 3647 1871 3657
rect 45 3637 1521 3647
rect 1541 3637 1621 3647
rect 45 3617 1511 3637
rect 1551 3627 1621 3637
rect 1681 3637 1741 3647
rect 1831 3637 1901 3647
rect 1981 3637 2451 3657
rect 2591 3647 3181 3657
rect 2601 3637 3191 3647
rect 1681 3627 1761 3637
rect 1851 3627 1911 3637
rect 1981 3627 2461 3637
rect 2621 3627 3201 3637
rect 3211 3627 3231 3637
rect 1561 3617 1631 3627
rect 1681 3617 1691 3627
rect 1711 3617 1781 3627
rect 45 3607 1501 3617
rect 1571 3607 1641 3617
rect 1731 3607 1791 3617
rect 1861 3607 1911 3627
rect 45 3597 1491 3607
rect 1591 3597 1671 3607
rect 45 3587 1501 3597
rect 1611 3587 1681 3597
rect 1741 3587 1801 3607
rect 1871 3597 1931 3607
rect 1901 3587 1941 3597
rect 1971 3587 2461 3627
rect 2631 3617 3231 3627
rect 2641 3607 2941 3617
rect 45 3577 1511 3587
rect 1521 3577 1561 3587
rect 1621 3577 1681 3587
rect 1751 3577 1811 3587
rect 1911 3582 2461 3587
rect 1911 3577 2321 3582
rect 2331 3577 2461 3582
rect 2651 3597 2941 3607
rect 2961 3597 3241 3617
rect 3391 3597 3411 3607
rect 2651 3587 3241 3597
rect 3351 3587 3371 3597
rect 2651 3577 3251 3587
rect 3291 3577 3301 3587
rect 3361 3577 3371 3587
rect 3381 3587 3411 3597
rect 3381 3577 3421 3587
rect 45 3567 1561 3577
rect 1631 3567 1681 3577
rect 1771 3567 1841 3577
rect 1921 3567 2301 3577
rect 2331 3567 2471 3577
rect 2651 3567 3321 3577
rect 3391 3567 3429 3577
rect 45 3547 1571 3567
rect 1631 3557 1691 3567
rect 1801 3557 1851 3567
rect 1931 3557 2291 3567
rect 2331 3557 2481 3567
rect 2651 3557 3011 3567
rect 3031 3557 3321 3567
rect 1641 3547 1731 3557
rect 1801 3547 1861 3557
rect 1931 3547 2491 3557
rect 2651 3547 3331 3557
rect 3411 3547 3429 3567
rect 45 3537 1581 3547
rect 1681 3537 1741 3547
rect 45 3527 1541 3537
rect 1571 3527 1621 3537
rect 1691 3527 1741 3537
rect 1811 3527 1861 3547
rect 1941 3537 2491 3547
rect 2641 3546 3345 3547
rect 3384 3546 3429 3547
rect 1931 3527 2481 3537
rect 2641 3527 3429 3546
rect 45 3497 1531 3527
rect 1571 3507 1631 3527
rect 1691 3517 1751 3527
rect 1831 3517 1851 3527
rect 1881 3517 1901 3527
rect 1931 3517 2471 3527
rect 2631 3517 2831 3527
rect 2841 3517 3321 3527
rect 1581 3497 1631 3507
rect 1701 3507 1751 3517
rect 1701 3497 1761 3507
rect 1871 3497 1911 3517
rect 1921 3497 2461 3517
rect 2621 3507 3331 3517
rect 3351 3507 3411 3527
rect 2611 3497 3421 3507
rect 45 3477 1541 3497
rect 1591 3495 1631 3497
rect 1591 3487 1620 3495
rect 1741 3487 1801 3497
rect 1611 3486 1620 3487
rect 1641 3486 1671 3487
rect 1611 3477 1621 3486
rect 1631 3477 1671 3486
rect 1751 3477 1801 3487
rect 1871 3477 2461 3497
rect 2481 3477 2501 3487
rect 2621 3477 3429 3497
rect 45 3467 1551 3477
rect 1631 3467 1681 3477
rect 1751 3467 1811 3477
rect 45 3447 1561 3467
rect 1631 3457 1691 3467
rect 1761 3457 1811 3467
rect 1641 3447 1691 3457
rect 1771 3447 1811 3457
rect 1891 3457 2511 3477
rect 2631 3457 3429 3477
rect 1891 3447 2521 3457
rect 2641 3447 3429 3457
rect 45 3427 1571 3447
rect 1641 3437 1710 3447
rect 1651 3427 1711 3437
rect 45 3377 1581 3427
rect 1677 3426 1741 3427
rect 1691 3417 1741 3426
rect 1821 3420 1861 3447
rect 1891 3437 2481 3447
rect 2491 3437 2511 3447
rect 1881 3420 2001 3437
rect 2011 3427 2431 3437
rect 1601 3397 1621 3407
rect 1701 3397 1751 3417
rect 1821 3407 2001 3420
rect 2021 3417 2431 3427
rect 2451 3427 2471 3437
rect 2651 3427 3429 3447
rect 2451 3417 2481 3427
rect 2671 3417 3429 3427
rect 1831 3405 2001 3407
rect 1831 3397 1851 3405
rect 1861 3397 2001 3405
rect 2031 3407 2481 3417
rect 2691 3407 3429 3417
rect 2031 3397 2491 3407
rect 2711 3397 2911 3407
rect 1601 3387 1631 3397
rect 1611 3384 1631 3387
rect 1711 3387 1761 3397
rect 1861 3387 2331 3397
rect 2341 3387 2501 3397
rect 2531 3387 2541 3396
rect 2721 3387 2911 3397
rect 2931 3387 3429 3407
rect 1611 3377 1623 3384
rect 1711 3377 1771 3387
rect 1861 3377 2501 3387
rect 2731 3377 2911 3387
rect 2921 3377 3429 3387
rect 45 3337 1591 3377
rect 1751 3367 1801 3377
rect 1861 3367 2511 3377
rect 2531 3367 2541 3377
rect 2741 3367 3429 3377
rect 1761 3357 1811 3367
rect 1861 3357 2021 3367
rect 2041 3357 2541 3367
rect 2751 3357 2941 3367
rect 1661 3347 1681 3357
rect 45 3327 1601 3337
rect 1651 3327 1691 3347
rect 1771 3337 1811 3357
rect 1851 3347 2021 3357
rect 2051 3347 2541 3357
rect 2761 3347 2931 3357
rect 1841 3337 2021 3347
rect 1781 3327 1811 3337
rect 1831 3327 2031 3337
rect 45 3307 1611 3327
rect 1661 3317 1691 3327
rect 1821 3317 2031 3327
rect 2061 3327 2551 3347
rect 2761 3337 2961 3347
rect 2971 3337 3429 3367
rect 2761 3327 3429 3337
rect 2061 3317 2381 3327
rect 2411 3317 2561 3327
rect 1681 3307 1691 3317
rect 1831 3307 1991 3317
rect 45 3267 1621 3307
rect 1931 3297 1991 3307
rect 2011 3307 2381 3317
rect 2421 3307 2561 3317
rect 2771 3307 3429 3327
rect 2011 3297 2341 3307
rect 1711 3287 1731 3297
rect 1941 3287 2001 3297
rect 2011 3287 2361 3297
rect 2431 3287 2461 3307
rect 2481 3297 2521 3307
rect 2531 3297 2571 3307
rect 2481 3287 2511 3297
rect 1711 3277 1751 3287
rect 1881 3277 1911 3287
rect 1941 3277 2361 3287
rect 1721 3267 1741 3277
rect 1871 3267 1921 3277
rect 45 3247 1631 3267
rect 1801 3257 1821 3267
rect 1791 3247 1821 3257
rect 1871 3257 1931 3267
rect 1941 3257 2041 3277
rect 2071 3267 2361 3277
rect 2381 3277 2391 3287
rect 2441 3277 2461 3287
rect 2491 3277 2511 3287
rect 2531 3287 2561 3297
rect 2641 3287 2651 3297
rect 2531 3277 2551 3287
rect 2381 3267 2401 3277
rect 2441 3267 2471 3277
rect 2481 3267 2511 3277
rect 1871 3247 1921 3257
rect 1951 3249 2041 3257
rect 2081 3257 2411 3267
rect 2441 3257 2521 3267
rect 2731 3257 2741 3267
rect 2781 3257 3429 3307
rect 1951 3247 2052 3249
rect 45 3227 1641 3247
rect 1781 3237 1811 3247
rect 1691 3227 1701 3237
rect 45 3197 1651 3227
rect 1891 3207 1911 3247
rect 1961 3237 2011 3247
rect 2031 3240 2052 3247
rect 1961 3227 2001 3237
rect 2031 3234 2058 3240
rect 2081 3237 2221 3257
rect 2040 3227 2058 3234
rect 2071 3227 2221 3237
rect 2231 3247 2411 3257
rect 2231 3237 2371 3247
rect 2231 3227 2241 3237
rect 2251 3227 2341 3237
rect 2351 3227 2361 3237
rect 1961 3207 2011 3227
rect 2040 3225 2361 3227
rect 2041 3207 2361 3225
rect 2381 3227 2421 3247
rect 2451 3237 2551 3257
rect 2591 3237 2611 3247
rect 2501 3227 2561 3237
rect 2381 3207 2431 3227
rect 2511 3217 2541 3227
rect 2601 3217 2611 3237
rect 2771 3227 3429 3257
rect 2781 3217 3429 3227
rect 2521 3207 2541 3217
rect 2781 3207 3041 3217
rect 1881 3197 1921 3207
rect 1951 3197 2231 3207
rect 45 3167 1661 3197
rect 1881 3187 1931 3197
rect 1941 3187 2231 3197
rect 1801 3177 1831 3187
rect 1881 3177 2061 3187
rect 2081 3177 2231 3187
rect 2241 3197 2331 3207
rect 2341 3197 2371 3207
rect 2241 3187 2371 3197
rect 2381 3197 2441 3207
rect 2381 3187 2451 3197
rect 2521 3187 2551 3207
rect 2781 3197 3001 3207
rect 3011 3197 3041 3207
rect 3051 3197 3429 3217
rect 2241 3177 2481 3187
rect 1721 3167 1731 3177
rect 45 3157 1671 3167
rect 1711 3157 1741 3167
rect 1801 3157 1841 3177
rect 1881 3167 2051 3177
rect 1881 3157 1931 3167
rect 1951 3157 2051 3167
rect 2081 3157 2481 3177
rect 2511 3157 2561 3187
rect 2601 3167 2611 3177
rect 2781 3167 3429 3197
rect 2601 3157 2621 3167
rect 2791 3157 3041 3167
rect 3051 3157 3429 3167
rect 45 3107 1681 3157
rect 1711 3137 1751 3157
rect 1811 3147 1831 3157
rect 1891 3137 1931 3157
rect 1961 3147 2021 3157
rect 2081 3147 2381 3157
rect 1721 3127 1751 3137
rect 1731 3107 1751 3127
rect 1901 3127 1931 3137
rect 1971 3127 2021 3147
rect 2071 3137 2381 3147
rect 2041 3127 2381 3137
rect 2391 3127 2471 3157
rect 2511 3147 2551 3157
rect 1901 3117 1941 3127
rect 1971 3117 2471 3127
rect 2521 3137 2551 3147
rect 2801 3137 3429 3157
rect 2521 3127 2541 3137
rect 2521 3117 2531 3127
rect 2811 3117 3429 3137
rect 1901 3107 1951 3117
rect 1971 3107 2481 3117
rect 45 3087 1691 3107
rect 1731 3097 1761 3107
rect 1901 3097 2381 3107
rect 2401 3097 2481 3107
rect 2681 3097 2691 3107
rect 2821 3097 3429 3117
rect 1731 3087 1771 3097
rect 1901 3087 1971 3097
rect 1981 3087 2381 3097
rect 45 3067 1701 3087
rect 45 3017 1711 3067
rect 1731 3057 1781 3087
rect 1831 3077 1851 3087
rect 1911 3077 1961 3087
rect 1981 3077 2061 3087
rect 1931 3067 1961 3077
rect 2001 3067 2061 3077
rect 2081 3077 2381 3087
rect 2411 3077 2491 3097
rect 2531 3087 2541 3097
rect 2601 3087 2621 3097
rect 2531 3077 2551 3087
rect 2601 3077 2631 3087
rect 2681 3077 2701 3097
rect 2831 3087 3429 3097
rect 2841 3077 3429 3087
rect 2081 3067 2491 3077
rect 2541 3067 2551 3077
rect 2611 3067 2631 3077
rect 2691 3067 2701 3077
rect 1951 3057 1971 3067
rect 2011 3057 2061 3067
rect 2091 3057 2501 3067
rect 2851 3057 3429 3077
rect 1741 3047 1781 3057
rect 1961 3047 1981 3057
rect 2021 3047 2071 3057
rect 2081 3047 2501 3057
rect 1751 3037 1781 3047
rect 1971 3037 2001 3047
rect 2021 3037 2501 3047
rect 1761 3017 1781 3037
rect 1981 3027 2011 3037
rect 2031 3027 2411 3037
rect 2421 3027 2511 3037
rect 1991 3017 2011 3027
rect 45 2997 1721 3017
rect 1761 3007 1791 3017
rect 1851 3007 1871 3017
rect 2001 3007 2021 3017
rect 2041 3007 2411 3027
rect 2431 3007 2511 3027
rect 45 2967 1731 2997
rect 1761 2967 1801 3007
rect 1851 2987 1881 3007
rect 1931 2997 1951 3007
rect 2001 2997 2031 3007
rect 2051 2997 2421 3007
rect 1941 2987 1961 2997
rect 2001 2987 2041 2997
rect 2051 2987 2081 2997
rect 2101 2987 2401 2997
rect 2431 2987 2521 3007
rect 2571 2997 2581 3007
rect 2631 2997 2651 3007
rect 2711 2997 2731 3017
rect 2861 3007 3429 3057
rect 2641 2987 2651 2997
rect 2011 2977 2081 2987
rect 2111 2977 2521 2987
rect 2871 2977 3429 3007
rect 2011 2967 2091 2977
rect 2111 2967 2531 2977
rect 45 2937 1741 2967
rect 1771 2957 1791 2967
rect 2021 2957 2421 2967
rect 2431 2957 2531 2967
rect 2881 2957 3429 2977
rect 2031 2947 2421 2957
rect 45 2907 1751 2937
rect 1881 2927 1901 2937
rect 1791 2917 1811 2927
rect 45 2897 1761 2907
rect 45 2857 1771 2897
rect 1781 2887 1821 2917
rect 1871 2907 1901 2927
rect 1961 2907 1981 2927
rect 2031 2917 2051 2947
rect 2061 2927 2421 2947
rect 2451 2947 2531 2957
rect 2891 2947 3429 2957
rect 2451 2937 2541 2947
rect 2901 2937 3429 2947
rect 2441 2927 2541 2937
rect 2591 2927 2611 2937
rect 2671 2927 2681 2937
rect 2031 2907 2061 2917
rect 2071 2907 2431 2927
rect 1881 2897 1891 2907
rect 2031 2897 2121 2907
rect 2031 2887 2131 2897
rect 2141 2887 2431 2907
rect 1801 2877 1811 2887
rect 2041 2867 2431 2887
rect 2451 2897 2551 2927
rect 2591 2917 2621 2927
rect 2741 2917 2761 2937
rect 2911 2927 3429 2937
rect 2931 2917 3429 2927
rect 2601 2907 2611 2917
rect 2941 2897 3429 2917
rect 2451 2877 2561 2897
rect 2951 2887 3429 2897
rect 45 2837 1781 2857
rect 1901 2847 1921 2857
rect 1811 2837 1831 2847
rect 45 2827 1791 2837
rect 1801 2827 1841 2837
rect 1891 2827 1931 2847
rect 1981 2837 2001 2847
rect 2041 2837 2061 2867
rect 2071 2857 2441 2867
rect 2481 2857 2561 2877
rect 2701 2857 2711 2867
rect 2961 2857 3429 2887
rect 2081 2847 2441 2857
rect 2081 2837 2431 2847
rect 2471 2837 2571 2857
rect 2611 2847 2631 2857
rect 2601 2837 2641 2847
rect 2691 2837 2721 2857
rect 2771 2837 2791 2857
rect 2841 2847 2851 2857
rect 2841 2837 2861 2847
rect 1991 2827 2011 2837
rect 45 2807 1841 2827
rect 1901 2817 1931 2827
rect 2041 2817 2071 2837
rect 2091 2827 2441 2837
rect 2081 2817 2451 2827
rect 2471 2817 2581 2837
rect 2611 2827 2641 2837
rect 2701 2827 2721 2837
rect 2971 2827 3429 2857
rect 2621 2817 2641 2827
rect 2041 2807 2451 2817
rect 2481 2807 2581 2817
rect 2961 2807 3429 2827
rect 45 2757 1811 2807
rect 2051 2787 2451 2807
rect 2491 2797 2581 2807
rect 2491 2787 2591 2797
rect 2061 2777 2081 2787
rect 2091 2777 2451 2787
rect 1911 2757 1941 2767
rect 45 2727 1861 2757
rect 1911 2737 1951 2757
rect 2011 2747 2021 2767
rect 2071 2757 2081 2777
rect 2111 2767 2301 2777
rect 2111 2757 2291 2767
rect 2311 2757 2461 2777
rect 2071 2747 2091 2757
rect 2121 2747 2291 2757
rect 2301 2747 2461 2757
rect 2501 2767 2591 2787
rect 2971 2777 3429 2807
rect 2711 2767 2731 2777
rect 2791 2767 2811 2777
rect 2971 2767 3181 2777
rect 3191 2767 3429 2777
rect 2071 2737 2101 2747
rect 2121 2737 2471 2747
rect 2501 2737 2601 2767
rect 2631 2737 2651 2767
rect 2701 2747 2741 2767
rect 2791 2757 2821 2767
rect 2861 2757 2881 2767
rect 2971 2757 3429 2767
rect 2801 2747 2811 2757
rect 2711 2737 2741 2747
rect 1921 2727 1951 2737
rect 2081 2727 2431 2737
rect 2451 2727 2461 2737
rect 2511 2727 2601 2737
rect 45 2717 1851 2727
rect 2091 2717 2111 2727
rect 2141 2717 2301 2727
rect 2311 2717 2471 2727
rect 2521 2717 2601 2727
rect 45 2697 1831 2717
rect 2151 2707 2301 2717
rect 2321 2707 2471 2717
rect 2511 2707 2611 2717
rect 2981 2707 3429 2757
rect 2151 2697 2411 2707
rect 2421 2697 2471 2707
rect 2521 2697 2611 2707
rect 45 2677 1841 2697
rect 1941 2677 1961 2687
rect 45 2667 1871 2677
rect 45 2637 1881 2667
rect 1931 2657 1971 2677
rect 2031 2667 2051 2687
rect 2151 2677 2481 2697
rect 2531 2687 2621 2697
rect 2521 2677 2621 2687
rect 2731 2677 2741 2687
rect 2811 2677 2831 2687
rect 2111 2667 2491 2677
rect 2031 2657 2061 2667
rect 2101 2657 2491 2667
rect 2531 2657 2621 2677
rect 2721 2667 2751 2677
rect 2801 2667 2841 2677
rect 2891 2667 2901 2687
rect 1941 2647 1971 2657
rect 2111 2647 2481 2657
rect 2531 2647 2631 2657
rect 2731 2647 2751 2667
rect 2811 2657 2841 2667
rect 2821 2647 2831 2657
rect 2121 2637 2491 2647
rect 45 2617 1871 2637
rect 2131 2627 2141 2637
rect 2151 2627 2491 2637
rect 2541 2627 2631 2647
rect 2151 2617 2501 2627
rect 2561 2617 2631 2627
rect 2991 2617 3429 2707
rect 45 2597 1861 2617
rect 2151 2607 2511 2617
rect 2561 2607 2641 2617
rect 2151 2597 2491 2607
rect 45 2587 1871 2597
rect 45 2497 1901 2587
rect 1951 2577 1991 2597
rect 2051 2577 2071 2597
rect 2121 2587 2141 2597
rect 2151 2587 2501 2597
rect 1961 2557 1991 2577
rect 2061 2567 2071 2577
rect 2111 2577 2501 2587
rect 2111 2567 2511 2577
rect 2561 2567 2651 2607
rect 2701 2577 2711 2597
rect 2761 2567 2771 2587
rect 2821 2567 2851 2597
rect 2911 2587 2921 2597
rect 2911 2577 2931 2587
rect 2921 2567 2931 2577
rect 2121 2547 2511 2567
rect 2151 2537 2521 2547
rect 2571 2537 2651 2567
rect 2831 2557 2841 2567
rect 3001 2557 3429 2617
rect 3011 2547 3429 2557
rect 3021 2537 3429 2547
rect 2151 2527 2531 2537
rect 2161 2517 2541 2527
rect 1981 2497 2011 2507
rect 45 2477 1921 2497
rect 1971 2487 2011 2497
rect 2071 2487 2091 2507
rect 2161 2497 2531 2517
rect 2561 2507 2651 2537
rect 3031 2517 3429 2537
rect 2701 2507 2721 2517
rect 2931 2507 2941 2517
rect 3041 2507 3429 2517
rect 45 2467 1931 2477
rect 1981 2467 2011 2487
rect 2081 2477 2091 2487
rect 2131 2477 2531 2497
rect 2551 2487 2661 2507
rect 2701 2487 2731 2507
rect 2841 2497 2861 2507
rect 2921 2497 2941 2507
rect 2781 2487 2791 2497
rect 2561 2477 2571 2487
rect 2141 2467 2531 2477
rect 2551 2467 2571 2477
rect 2581 2467 2661 2487
rect 2841 2477 2871 2497
rect 2921 2487 2951 2497
rect 3031 2487 3429 2507
rect 2931 2477 2941 2487
rect 3041 2467 3429 2487
rect 45 2427 1921 2467
rect 2141 2457 2661 2467
rect 3051 2457 3429 2467
rect 2151 2447 2661 2457
rect 2161 2437 2671 2447
rect 3061 2437 3429 2457
rect 2171 2427 2671 2437
rect 45 2407 1931 2427
rect 2171 2417 2661 2427
rect 2711 2417 2731 2427
rect 2941 2417 2951 2427
rect 3011 2417 3021 2427
rect 3071 2417 3429 2437
rect 2001 2407 2031 2417
rect 2091 2407 2111 2417
rect 45 2377 1941 2407
rect 1991 2397 2041 2407
rect 2001 2387 2041 2397
rect 2091 2387 2121 2407
rect 2001 2377 2031 2387
rect 2161 2377 2671 2417
rect 2711 2387 2741 2417
rect 2791 2397 2811 2417
rect 2861 2397 2881 2417
rect 2931 2397 2961 2417
rect 2801 2387 2811 2397
rect 2871 2387 2891 2397
rect 2941 2387 2961 2397
rect 3011 2387 3031 2417
rect 3061 2407 3429 2417
rect 3071 2377 3429 2407
rect 45 2327 1951 2377
rect 2171 2367 2681 2377
rect 2171 2357 2671 2367
rect 2181 2347 2671 2357
rect 45 2297 1961 2327
rect 2021 2317 2041 2327
rect 2111 2317 2131 2327
rect 2021 2297 2051 2317
rect 2111 2307 2141 2317
rect 2181 2307 2681 2347
rect 3081 2337 3429 2377
rect 2721 2327 2731 2337
rect 2791 2327 2811 2337
rect 2871 2327 2881 2337
rect 2711 2307 2741 2327
rect 2121 2297 2131 2307
rect 45 2257 1971 2297
rect 2031 2287 2051 2297
rect 2181 2287 2571 2307
rect 2581 2287 2681 2307
rect 2721 2297 2741 2307
rect 2791 2307 2821 2327
rect 2791 2297 2811 2307
rect 2861 2297 2891 2327
rect 2941 2317 2961 2327
rect 3011 2317 3031 2327
rect 2931 2307 2961 2317
rect 3001 2307 3031 2317
rect 2941 2297 2961 2307
rect 3011 2297 3031 2307
rect 3071 2317 3321 2337
rect 3341 2327 3429 2337
rect 3331 2317 3429 2327
rect 2871 2287 2881 2297
rect 3071 2287 3429 2317
rect 2181 2277 2681 2287
rect 3071 2277 3321 2287
rect 2191 2267 2681 2277
rect 3081 2267 3311 2277
rect 3341 2267 3429 2287
rect 2191 2257 2581 2267
rect 45 2237 1981 2257
rect 2191 2247 2571 2257
rect 2591 2247 2691 2267
rect 45 2197 1991 2237
rect 2051 2227 2071 2237
rect 2131 2227 2151 2237
rect 2051 2217 2081 2227
rect 2141 2217 2151 2227
rect 2191 2235 2691 2247
rect 2701 2235 2741 2237
rect 2061 2207 2071 2217
rect 2191 2207 2741 2235
rect 2191 2205 2730 2207
rect 2191 2197 2709 2205
rect 2791 2197 2811 2237
rect 2861 2227 2881 2247
rect 2941 2237 2951 2247
rect 3011 2237 3021 2247
rect 2851 2217 2881 2227
rect 2861 2197 2881 2217
rect 2931 2227 2951 2237
rect 2931 2217 2961 2227
rect 2931 2197 2951 2217
rect 3001 2207 3031 2237
rect 3071 2227 3429 2267
rect 3061 2217 3341 2227
rect 3351 2217 3429 2227
rect 3001 2197 3021 2207
rect 3061 2197 3429 2217
rect 45 2167 2001 2197
rect 2201 2187 2561 2197
rect 2571 2190 2709 2197
rect 2571 2187 2701 2190
rect 2201 2177 2701 2187
rect 45 2137 2011 2167
rect 2071 2147 2091 2157
rect 2211 2147 2701 2177
rect 3071 2187 3429 2197
rect 3071 2157 3121 2187
rect 3131 2157 3429 2187
rect 2061 2137 2091 2147
rect 45 2117 2021 2137
rect 2071 2117 2091 2137
rect 2151 2137 2161 2147
rect 2211 2137 2721 2147
rect 2151 2117 2171 2137
rect 2211 2127 2741 2137
rect 2791 2127 2811 2147
rect 2861 2127 2881 2147
rect 2931 2127 2951 2147
rect 2211 2117 2731 2127
rect 2801 2117 2811 2127
rect 2871 2117 2881 2127
rect 2941 2117 2951 2127
rect 3001 2137 3021 2147
rect 3061 2137 3429 2157
rect 3001 2117 3031 2137
rect 3051 2127 3429 2137
rect 3041 2117 3429 2127
rect 45 2107 2011 2117
rect 2221 2107 2701 2117
rect 3011 2107 3021 2117
rect 3051 2107 3429 2117
rect 45 2077 2021 2107
rect 2221 2097 2711 2107
rect 2231 2077 2711 2097
rect 3061 2087 3429 2107
rect 45 2047 2031 2077
rect 2241 2067 2681 2077
rect 2691 2067 2721 2077
rect 3071 2067 3111 2087
rect 3131 2067 3429 2087
rect 45 2007 2041 2047
rect 2081 2027 2101 2057
rect 2151 2047 2171 2057
rect 2231 2047 2681 2067
rect 2701 2047 2711 2067
rect 2151 2027 2181 2047
rect 2221 2037 2721 2047
rect 2221 2027 2401 2037
rect 2411 2027 2421 2037
rect 2431 2027 2721 2037
rect 2741 2027 2761 2057
rect 2811 2047 2831 2057
rect 2811 2037 2841 2047
rect 2881 2037 2901 2057
rect 2821 2027 2841 2037
rect 2891 2027 2911 2037
rect 2951 2027 2971 2057
rect 3011 2047 3041 2057
rect 3061 2047 3429 2067
rect 3011 2037 3429 2047
rect 3011 2027 3041 2037
rect 2161 2017 2171 2027
rect 2221 2017 2721 2027
rect 2961 2017 2971 2027
rect 3021 2017 3041 2027
rect 3051 2017 3429 2037
rect 45 1987 2051 2007
rect 2231 1997 2731 2017
rect 3021 2007 3031 2017
rect 45 1947 2061 1987
rect 2231 1977 2721 1997
rect 3061 1987 3429 2017
rect 3061 1977 3101 1987
rect 3111 1977 3429 1987
rect 2231 1967 2731 1977
rect 2821 1967 2831 1977
rect 3031 1967 3041 1977
rect 3061 1967 3429 1977
rect 45 1927 2071 1947
rect 2091 1937 2111 1967
rect 2231 1957 2761 1967
rect 2161 1927 2181 1957
rect 2221 1947 2771 1957
rect 2221 1937 2761 1947
rect 2811 1937 2841 1967
rect 2891 1957 2911 1967
rect 2971 1957 2981 1967
rect 2891 1937 2921 1957
rect 2961 1937 2981 1957
rect 3021 1937 3429 1967
rect 2221 1927 2731 1937
rect 2891 1927 2911 1937
rect 45 1897 2081 1927
rect 2231 1917 2731 1927
rect 3031 1917 3429 1937
rect 2241 1907 2741 1917
rect 3041 1907 3051 1917
rect 2271 1897 2741 1907
rect 3071 1897 3429 1917
rect 45 1877 2091 1897
rect 45 1857 2111 1877
rect 2281 1867 2741 1897
rect 3041 1887 3051 1897
rect 3041 1877 3061 1887
rect 3081 1877 3429 1897
rect 45 1847 2121 1857
rect 2171 1847 2181 1867
rect 2241 1857 2261 1867
rect 2271 1857 2401 1867
rect 2411 1857 2771 1867
rect 2231 1847 2771 1857
rect 2821 1847 2841 1877
rect 2891 1867 2911 1877
rect 2971 1867 2991 1877
rect 2891 1847 2921 1867
rect 2961 1847 2991 1867
rect 45 1807 2111 1847
rect 2171 1837 2191 1847
rect 2231 1837 2741 1847
rect 2901 1837 2911 1847
rect 2971 1837 2991 1847
rect 3041 1837 3429 1877
rect 2241 1827 2251 1837
rect 2271 1827 2741 1837
rect 45 1787 2121 1807
rect 2291 1787 2741 1827
rect 3041 1807 3071 1837
rect 3081 1827 3429 1837
rect 3051 1797 3071 1807
rect 3091 1797 3429 1827
rect 45 1757 2131 1787
rect 2181 1767 2191 1777
rect 2291 1767 2751 1787
rect 2911 1777 2921 1787
rect 2981 1777 2991 1787
rect 45 1727 2141 1757
rect 2181 1747 2201 1767
rect 2251 1757 2461 1767
rect 2471 1757 2751 1767
rect 2791 1757 2801 1777
rect 2841 1767 2861 1777
rect 2851 1757 2861 1767
rect 2911 1757 2931 1777
rect 2971 1767 3001 1777
rect 2251 1737 2741 1757
rect 2981 1747 3001 1767
rect 3041 1747 3429 1797
rect 3041 1737 3101 1747
rect 45 1697 2151 1727
rect 2291 1717 2751 1737
rect 2301 1707 2751 1717
rect 3051 1707 3091 1737
rect 45 1677 2161 1697
rect 2301 1687 2761 1707
rect 3051 1697 3101 1707
rect 3111 1697 3429 1747
rect 2261 1677 2271 1687
rect 2291 1677 2761 1687
rect 45 1667 2171 1677
rect 45 1577 2161 1667
rect 2191 1647 2211 1677
rect 2251 1667 2431 1677
rect 2441 1667 2761 1677
rect 2791 1687 2811 1697
rect 2791 1667 2821 1687
rect 2861 1677 2881 1697
rect 2991 1687 3001 1697
rect 2871 1667 2881 1677
rect 2921 1667 2941 1687
rect 2251 1657 2411 1667
rect 2501 1657 2531 1667
rect 2551 1657 2761 1667
rect 2991 1657 3011 1687
rect 3041 1657 3429 1697
rect 2261 1647 2401 1657
rect 2671 1647 2771 1657
rect 3051 1647 3429 1657
rect 2291 1637 2381 1647
rect 2301 1627 2371 1637
rect 2201 1577 2211 1587
rect 2301 1577 2381 1627
rect 3051 1617 3111 1647
rect 3121 1617 3429 1647
rect 2811 1587 2821 1607
rect 2871 1577 2891 1607
rect 2941 1597 2951 1607
rect 2931 1587 2961 1597
rect 2941 1577 2961 1587
rect 45 1567 2171 1577
rect 45 1527 2161 1567
rect 2201 1557 2221 1577
rect 2261 1567 2281 1577
rect 2291 1567 2431 1577
rect 2451 1567 2601 1577
rect 2871 1567 2881 1577
rect 2941 1567 2951 1577
rect 3001 1567 3021 1597
rect 3051 1587 3429 1617
rect 3041 1567 3429 1587
rect 2261 1547 2781 1567
rect 3051 1557 3429 1567
rect 2301 1537 2591 1547
rect 2601 1537 2781 1547
rect 2301 1527 2541 1537
rect 2561 1527 2591 1537
rect 2611 1527 2651 1537
rect 45 1487 2171 1527
rect 2311 1497 2541 1527
rect 2551 1517 2601 1527
rect 2611 1517 2641 1527
rect 2661 1517 2781 1537
rect 3061 1537 3429 1557
rect 3061 1527 3111 1537
rect 3131 1527 3429 1537
rect 2551 1507 2791 1517
rect 3061 1507 3429 1527
rect 2551 1497 2771 1507
rect 2831 1497 2841 1507
rect 2211 1487 2221 1497
rect 45 1407 2181 1487
rect 2201 1467 2221 1487
rect 2271 1487 2291 1497
rect 2311 1487 2771 1497
rect 2891 1487 2901 1507
rect 2951 1497 2961 1507
rect 2951 1487 2971 1497
rect 2271 1477 2651 1487
rect 2661 1477 2791 1487
rect 2951 1477 2961 1487
rect 3011 1477 3429 1507
rect 2271 1467 2771 1477
rect 3021 1467 3041 1477
rect 2271 1457 2281 1467
rect 2311 1437 2791 1467
rect 3061 1457 3429 1477
rect 2321 1417 2801 1437
rect 2321 1407 2791 1417
rect 45 1397 2191 1407
rect 2321 1397 2811 1407
rect 2841 1397 2861 1427
rect 2901 1417 2911 1427
rect 3031 1417 3051 1427
rect 3071 1417 3429 1457
rect 2901 1397 2921 1417
rect 45 1327 2201 1397
rect 2211 1367 2231 1397
rect 2281 1387 2791 1397
rect 2911 1387 2921 1397
rect 2961 1387 2981 1417
rect 2271 1377 2791 1387
rect 2801 1377 2811 1387
rect 3021 1377 3429 1417
rect 2281 1367 2821 1377
rect 2281 1357 2831 1367
rect 2311 1347 2821 1357
rect 2321 1337 2821 1347
rect 3031 1337 3051 1377
rect 2321 1327 2831 1337
rect 2841 1327 2861 1337
rect 2911 1327 2921 1337
rect 3021 1327 3051 1337
rect 3071 1327 3429 1377
rect 45 1307 2211 1327
rect 2321 1307 2861 1327
rect 2901 1307 2921 1327
rect 2971 1317 2981 1327
rect 45 1297 2221 1307
rect 2281 1297 2861 1307
rect 2911 1297 2921 1307
rect 2961 1297 2981 1317
rect 45 1267 2231 1297
rect 2281 1287 2841 1297
rect 3021 1287 3429 1327
rect 2281 1277 2851 1287
rect 45 1237 2221 1267
rect 2291 1257 2851 1277
rect 2331 1247 2851 1257
rect 2331 1237 2611 1247
rect 2631 1237 2851 1247
rect 3021 1237 3051 1287
rect 3061 1277 3429 1287
rect 3071 1237 3429 1277
rect 45 1207 2231 1237
rect 2331 1227 2561 1237
rect 2581 1227 2641 1237
rect 2651 1227 2861 1237
rect 2911 1227 2921 1237
rect 2331 1207 2541 1227
rect 2571 1217 2641 1227
rect 2561 1207 2651 1217
rect 2661 1207 2861 1227
rect 2901 1207 2921 1227
rect 2971 1217 2981 1237
rect 3021 1217 3429 1237
rect 2961 1207 2981 1217
rect 45 1117 2241 1207
rect 2291 1197 2541 1207
rect 2281 1177 2541 1197
rect 2551 1187 2861 1207
rect 2911 1197 2921 1207
rect 2971 1197 2981 1207
rect 3011 1197 3429 1217
rect 3021 1187 3429 1197
rect 2561 1177 2851 1187
rect 2291 1167 2851 1177
rect 2301 1157 2321 1167
rect 2331 1157 2851 1167
rect 3021 1157 3051 1187
rect 3061 1177 3429 1187
rect 2331 1147 2861 1157
rect 3011 1147 3051 1157
rect 3071 1147 3429 1177
rect 2291 1117 2321 1127
rect 2341 1117 2861 1147
rect 2901 1137 2921 1147
rect 2891 1117 2921 1137
rect 45 1057 2251 1117
rect 2281 1077 2861 1117
rect 2901 1107 2921 1117
rect 2961 1107 2981 1137
rect 3011 1117 3429 1147
rect 3001 1107 3429 1117
rect 2291 1067 2861 1077
rect 45 1027 2261 1057
rect 2291 1047 2311 1067
rect 2301 1037 2311 1047
rect 2331 1037 2861 1067
rect 3011 1097 3429 1107
rect 3011 1087 3051 1097
rect 3011 1067 3041 1087
rect 3011 1057 3051 1067
rect 3061 1057 3429 1097
rect 2891 1047 2911 1057
rect 2301 1027 2321 1037
rect 2331 1027 2871 1037
rect 45 977 2271 1027
rect 2291 1017 2871 1027
rect 2881 1027 2921 1047
rect 2961 1037 2981 1047
rect 3001 1037 3429 1057
rect 2881 1017 2911 1027
rect 2961 1017 3429 1037
rect 2291 997 2861 1017
rect 2891 1007 2911 1017
rect 2971 1007 3429 1017
rect 3001 997 3429 1007
rect 2301 987 2861 997
rect 2311 977 2861 987
rect 45 937 2281 977
rect 2321 967 2331 977
rect 2341 967 2871 977
rect 3011 967 3041 997
rect 3051 967 3429 997
rect 2341 957 2911 967
rect 2351 947 2911 957
rect 2321 937 2331 947
rect 2341 937 2911 947
rect 2961 957 2991 967
rect 3001 957 3429 967
rect 2961 937 3429 957
rect 45 917 2291 937
rect 2311 927 2911 937
rect 2311 917 2901 927
rect 2951 917 3429 937
rect 45 887 2871 917
rect 45 877 2341 887
rect 45 857 2311 877
rect 2321 867 2341 877
rect 2331 857 2341 867
rect 45 847 2341 857
rect 2351 877 2871 887
rect 2961 877 2981 917
rect 2351 867 2891 877
rect 2951 867 2981 877
rect 3001 897 3429 917
rect 3001 877 3041 897
rect 3051 877 3429 897
rect 2351 847 2901 867
rect 2951 857 2991 867
rect 3001 857 3429 877
rect 45 837 2901 847
rect 45 827 2891 837
rect 45 797 2871 827
rect 2941 817 3429 857
rect 45 787 2341 797
rect 2351 787 2881 797
rect 2941 787 2981 817
rect 45 777 2331 787
rect 2361 777 2881 787
rect 2931 777 2981 787
rect 3001 807 3429 817
rect 3001 787 3041 807
rect 3051 787 3429 807
rect 3001 777 3429 787
rect 45 747 2341 777
rect 2361 767 2891 777
rect 2921 767 2981 777
rect 2991 767 3429 777
rect 2361 747 2881 767
rect 2921 757 3429 767
rect 2911 747 3429 757
rect 45 737 2881 747
rect 2921 737 3429 747
rect 45 677 2871 737
rect 2921 727 2981 737
rect 2921 687 2971 727
rect 2991 707 3429 737
rect 3001 697 3429 707
rect 2901 677 2971 687
rect 2991 677 3429 697
rect 45 667 2881 677
rect 2891 667 3429 677
rect 45 657 3429 667
rect 45 647 2881 657
rect 2891 647 3429 657
rect 45 627 2871 647
rect 2911 637 3429 647
rect 2911 627 2961 637
rect 2981 627 3429 637
rect 45 597 2881 627
rect 2921 617 2961 627
rect 2911 597 2961 617
rect 2991 597 3429 627
rect 45 587 2891 597
rect 2901 587 2961 597
rect 2981 587 3429 597
rect 45 557 3429 587
rect 45 497 2881 557
rect 2901 547 3429 557
rect 2901 537 2961 547
rect 2901 507 2951 537
rect 2891 497 2951 507
rect 2981 497 3429 547
rect 45 457 3429 497
rect 45 447 2951 457
rect 45 417 2881 447
rect 2891 417 2941 447
rect 45 407 2941 417
rect 2971 407 3429 457
rect 45 397 2951 407
rect 2961 397 3429 407
rect 45 367 3429 397
rect 45 357 2941 367
rect 2951 357 3429 367
rect 45 317 2931 357
rect 2961 317 3429 357
rect 45 267 3429 317
rect 45 257 2931 267
rect 2941 257 3429 267
rect 45 227 2921 257
rect 2951 237 3429 257
rect 2941 227 3429 237
rect 45 167 3429 227
rect 45 147 2911 167
rect 2931 147 3429 167
rect 45 87 3429 147
use evan-threshold  evan-threshold_0
timestamp 1419145638
transform 1 0 2770 0 1 93
box 515 -15 7873 7185
<< end >>
