magic
tech scmos
timestamp 1418688738
<< electrode >>
rect 96 -170 102 -163
rect 96 -201 102 -194
<< electrodecontact >>
rect 97 -168 101 -164
rect 97 -200 101 -196
<< ntransistor >>
rect 27 -156 33 -36
rect 39 -156 45 -36
rect 51 -156 57 -36
rect 63 -156 69 -36
rect 83 -276 89 -36
rect 101 -156 107 -36
rect 121 -156 127 -36
rect 133 -156 139 -36
rect 145 -156 151 -36
rect 157 -156 163 -36
<< ptransistor >>
rect 27 -24 33 96
rect 39 -24 45 96
rect 51 -24 57 96
rect 63 -24 69 96
rect 83 -24 89 96
rect 101 -24 107 96
rect 121 -24 127 96
rect 133 -24 139 96
rect 145 -24 151 96
rect 157 -24 163 96
<< ndiffusion >>
rect 24 -38 27 -36
rect 26 -42 27 -38
rect 24 -156 27 -42
rect 33 -44 39 -36
rect 33 -48 34 -44
rect 38 -48 39 -44
rect 33 -156 39 -48
rect 45 -37 51 -36
rect 45 -41 46 -37
rect 50 -41 51 -37
rect 45 -156 51 -41
rect 57 -44 63 -36
rect 57 -48 58 -44
rect 62 -48 63 -44
rect 57 -156 63 -48
rect 69 -43 72 -36
rect 82 -40 83 -36
rect 69 -47 70 -43
rect 69 -156 72 -47
rect 80 -276 83 -40
rect 89 -196 92 -36
rect 98 -43 101 -36
rect 100 -47 101 -43
rect 98 -152 101 -47
rect 100 -156 101 -152
rect 107 -40 108 -36
rect 120 -40 121 -36
rect 107 -152 110 -40
rect 107 -156 108 -152
rect 118 -156 121 -40
rect 127 -156 133 -36
rect 139 -156 145 -36
rect 151 -43 157 -36
rect 151 -47 152 -43
rect 156 -47 157 -43
rect 151 -156 157 -47
rect 163 -38 166 -36
rect 163 -42 164 -38
rect 163 -156 166 -42
rect 89 -200 90 -196
rect 89 -276 92 -200
<< pdiffusion >>
rect 24 -18 27 96
rect 26 -22 27 -18
rect 24 -24 27 -22
rect 33 -13 39 96
rect 33 -17 34 -13
rect 38 -17 39 -13
rect 33 -24 39 -17
rect 45 -24 51 96
rect 57 -24 63 96
rect 69 -20 72 96
rect 82 92 83 96
rect 80 -20 83 92
rect 69 -24 70 -20
rect 82 -24 83 -20
rect 89 -13 92 96
rect 98 -13 101 96
rect 89 -17 90 -13
rect 100 -17 101 -13
rect 89 -24 92 -17
rect 98 -24 101 -17
rect 107 -20 110 96
rect 118 -13 121 96
rect 120 -17 121 -13
rect 107 -24 108 -20
rect 118 -24 121 -17
rect 127 -12 133 96
rect 127 -16 128 -12
rect 132 -16 133 -12
rect 127 -24 133 -16
rect 139 -19 145 96
rect 139 -23 140 -19
rect 144 -23 145 -19
rect 139 -24 145 -23
rect 151 -12 157 96
rect 151 -16 152 -12
rect 156 -16 157 -12
rect 151 -24 157 -16
rect 163 -18 166 96
rect 163 -22 164 -18
rect 163 -24 166 -22
<< ndcontact >>
rect 22 -42 26 -38
rect 34 -48 38 -44
rect 46 -41 50 -37
rect 58 -48 62 -44
rect 78 -40 82 -36
rect 70 -47 74 -43
rect 96 -47 100 -43
rect 96 -156 100 -152
rect 108 -40 112 -36
rect 116 -40 120 -36
rect 108 -156 112 -152
rect 152 -47 156 -43
rect 164 -42 168 -38
rect 90 -200 94 -196
<< pdcontact >>
rect 22 -22 26 -18
rect 34 -17 38 -13
rect 78 92 82 96
rect 70 -24 74 -20
rect 78 -24 82 -20
rect 90 -17 100 -13
rect 116 -17 120 -13
rect 108 -24 112 -20
rect 128 -16 132 -12
rect 140 -23 144 -19
rect 152 -16 156 -12
rect 164 -22 168 -18
<< polysilicon >>
rect 27 97 64 99
rect 68 97 69 99
rect 27 96 33 97
rect 39 96 45 97
rect 51 96 57 97
rect 63 96 69 97
rect 83 96 89 98
rect 101 96 107 98
rect 121 96 127 99
rect 133 96 139 99
rect 145 96 151 99
rect 157 96 163 99
rect 27 -26 33 -24
rect 39 -26 45 -24
rect 51 -26 57 -24
rect 63 -26 69 -24
rect 83 -25 89 -24
rect 101 -25 107 -24
rect 83 -27 84 -25
rect 88 -27 107 -25
rect 121 -25 127 -24
rect 133 -25 139 -24
rect 145 -25 151 -24
rect 121 -27 122 -25
rect 126 -27 140 -25
rect 144 -27 151 -25
rect 157 -25 163 -24
rect 157 -26 158 -25
rect 162 -26 163 -25
rect 27 -35 28 -34
rect 32 -35 33 -34
rect 27 -36 33 -35
rect 39 -35 46 -33
rect 50 -35 64 -33
rect 68 -35 69 -34
rect 39 -36 45 -35
rect 51 -36 57 -35
rect 63 -36 69 -35
rect 83 -35 102 -33
rect 106 -35 107 -33
rect 83 -36 89 -35
rect 101 -36 107 -35
rect 121 -36 127 -34
rect 133 -36 139 -34
rect 145 -36 151 -34
rect 157 -36 163 -34
rect 27 -158 33 -156
rect 39 -158 45 -156
rect 51 -158 57 -156
rect 63 -158 69 -156
rect 101 -158 107 -156
rect 121 -157 127 -156
rect 133 -157 139 -156
rect 145 -157 151 -156
rect 157 -157 163 -156
rect 121 -159 122 -157
rect 126 -159 163 -157
rect 83 -278 89 -276
<< polycontact >>
rect 64 97 68 101
rect 84 -29 88 -25
rect 122 -29 126 -25
rect 140 -29 144 -25
rect 158 -29 162 -25
rect 28 -35 32 -31
rect 46 -35 50 -31
rect 64 -35 68 -31
rect 102 -35 106 -31
rect 122 -161 126 -157
<< metal1 >>
rect 68 97 82 101
rect 78 96 82 97
rect 38 -17 90 -13
rect 100 -17 116 -13
rect 132 -16 152 -12
rect 22 -31 26 -22
rect 70 -31 74 -24
rect 22 -35 28 -31
rect 68 -35 74 -31
rect 78 -25 82 -24
rect 78 -29 84 -25
rect 22 -38 26 -35
rect 46 -37 50 -35
rect 78 -36 82 -29
rect 108 -31 112 -24
rect 140 -25 144 -23
rect 164 -25 168 -22
rect 106 -35 112 -31
rect 108 -36 112 -35
rect 116 -29 122 -25
rect 162 -29 168 -25
rect 116 -36 120 -29
rect 164 -38 168 -29
rect 38 -48 58 -44
rect 74 -47 96 -43
rect 100 -47 152 -43
rect 96 -164 100 -156
rect 108 -157 112 -156
rect 108 -161 122 -157
rect 96 -168 97 -164
rect 94 -200 97 -196
<< high_resist >>
rect 94 -194 96 -170
rect 102 -194 104 -170
<< poly2_high_resist >>
rect 96 -194 102 -170
<< labels >>
rlabel polysilicon 63 97 69 99 5 Vbp
rlabel metal1 22 -35 26 -31 3 Vcn
rlabel metal1 78 -36 82 -24 1 Vbp
rlabel metal1 108 -36 112 -24 1 Vbn
rlabel metal1 164 -29 168 -25 7 Vcp
rlabel polysilicon 121 -159 127 -157 1 Vbn
rlabel pdcontact 116 -17 120 -13 1 Vdd
rlabel pdcontact 34 -17 38 -13 1 Vdd
rlabel ndcontact 152 -47 156 -43 1 Gnd
rlabel ndcontact 70 -47 74 -43 1 Gnd
<< end >>
