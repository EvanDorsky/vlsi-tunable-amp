magic
tech scmos
timestamp 1418852285
<< nwell >>
rect 58 0 62 3
rect 43 -4 86 0
rect 142 0 146 1
rect 129 -4 172 0
rect 0 -136 2 -4
rect 58 -5 62 -4
rect 153 -5 157 -4
rect 231 -119 1624 137
<< pwell >>
rect 0 -4 43 3
rect 86 -4 129 3
rect 0 -388 2 -136
rect 231 -373 1449 -119
<< electrodecontact >>
rect 1000 60 1004 212
rect 852 -107 856 43
<< electrodecap >>
rect 850 58 1006 214
rect 850 -111 1006 45
<< ntransistor >>
rect 243 -367 249 -127
rect 255 -367 261 -127
rect 267 -367 273 -127
rect 279 -367 285 -127
rect 291 -367 297 -127
rect 303 -367 309 -127
rect 315 -367 321 -127
rect 327 -367 333 -127
rect 339 -367 345 -127
rect 351 -367 357 -127
rect 363 -367 369 -127
rect 375 -367 381 -127
rect 387 -367 393 -127
rect 399 -367 405 -127
rect 411 -367 417 -127
rect 423 -367 429 -127
rect 435 -367 441 -127
rect 447 -367 453 -127
rect 459 -367 465 -127
rect 471 -367 477 -127
rect 483 -367 489 -127
rect 495 -367 501 -127
rect 507 -367 513 -127
rect 519 -367 525 -127
rect 531 -367 537 -127
rect 543 -367 549 -127
rect 555 -367 561 -127
rect 567 -367 573 -127
rect 579 -367 585 -127
rect 591 -367 597 -127
rect 603 -367 609 -127
rect 615 -367 621 -127
rect 627 -367 633 -127
rect 639 -367 645 -127
rect 651 -367 657 -127
rect 663 -367 669 -127
rect 675 -367 681 -127
rect 687 -367 693 -127
rect 699 -367 705 -127
rect 711 -367 717 -127
rect 723 -367 729 -127
rect 735 -367 741 -127
rect 747 -367 753 -127
rect 759 -367 765 -127
rect 771 -367 777 -127
rect 783 -367 789 -127
rect 795 -367 801 -127
rect 807 -367 813 -127
rect 819 -367 825 -127
rect 831 -367 837 -127
rect 843 -367 849 -127
rect 855 -367 861 -127
rect 867 -367 873 -127
rect 879 -367 885 -127
rect 891 -367 897 -127
rect 903 -367 909 -127
rect 915 -367 921 -127
rect 927 -367 933 -127
rect 939 -367 945 -127
rect 951 -367 957 -127
rect 963 -367 969 -127
rect 975 -367 981 -127
rect 987 -367 993 -127
rect 999 -367 1005 -127
rect 1011 -367 1017 -127
rect 1023 -367 1029 -127
rect 1035 -367 1041 -127
rect 1047 -367 1053 -127
rect 1059 -367 1065 -127
rect 1071 -367 1077 -127
rect 1083 -367 1089 -127
rect 1095 -367 1101 -127
rect 1107 -367 1113 -127
rect 1119 -367 1125 -127
rect 1131 -367 1137 -127
rect 1143 -367 1149 -127
rect 1155 -367 1161 -127
rect 1167 -367 1173 -127
rect 1179 -367 1185 -127
rect 1191 -367 1197 -127
rect 1203 -367 1209 -127
rect 1215 -367 1221 -127
rect 1227 -367 1233 -127
rect 1239 -367 1245 -127
rect 1251 -367 1257 -127
rect 1263 -367 1269 -127
rect 1275 -367 1281 -127
rect 1287 -367 1293 -127
rect 1299 -367 1305 -127
rect 1311 -367 1317 -127
rect 1323 -367 1329 -127
rect 1335 -367 1341 -127
rect 1347 -367 1353 -127
rect 1359 -367 1365 -127
rect 1371 -367 1377 -127
rect 1383 -367 1389 -127
rect 1395 -367 1401 -127
rect 1407 -367 1413 -127
rect 1419 -367 1425 -127
rect 1431 -367 1437 -127
<< ptransistor >>
rect 243 -109 249 131
rect 255 -109 261 131
rect 267 -109 273 131
rect 279 -109 285 131
rect 291 -109 297 131
rect 303 -109 309 131
rect 315 -109 321 131
rect 327 -109 333 131
rect 339 -109 345 131
rect 351 -109 357 131
rect 363 -109 369 131
rect 375 -109 381 131
rect 387 -109 393 131
rect 399 -109 405 131
rect 411 -109 417 131
rect 423 -109 429 131
rect 435 -109 441 131
rect 447 -109 453 131
rect 459 -109 465 131
rect 471 -109 477 131
rect 483 -109 489 131
rect 495 -109 501 131
rect 507 -109 513 131
rect 519 -109 525 131
rect 531 -109 537 131
rect 543 -109 549 131
rect 555 -109 561 131
rect 567 -109 573 131
rect 579 -109 585 131
rect 591 -109 597 131
rect 603 -109 609 131
rect 615 -109 621 131
rect 627 -109 633 131
rect 639 -109 645 131
rect 651 -109 657 131
rect 663 -109 669 131
rect 675 -109 681 131
rect 687 -109 693 131
rect 699 -109 705 131
rect 711 -109 717 131
rect 723 -109 729 131
rect 735 -109 741 131
rect 747 -109 753 131
rect 759 -109 765 131
rect 771 -109 777 131
rect 783 -109 789 131
rect 795 -109 801 131
rect 807 -109 813 131
rect 819 -109 825 131
rect 831 -109 837 131
rect 1018 -109 1024 131
rect 1030 -109 1036 131
rect 1042 -109 1048 131
rect 1054 -109 1060 131
rect 1066 -109 1072 131
rect 1078 -109 1084 131
rect 1090 -109 1096 131
rect 1102 -109 1108 131
rect 1114 -109 1120 131
rect 1126 -109 1132 131
rect 1138 -109 1144 131
rect 1150 -109 1156 131
rect 1162 -109 1168 131
rect 1174 -109 1180 131
rect 1186 -109 1192 131
rect 1198 -109 1204 131
rect 1210 -109 1216 131
rect 1222 -109 1228 131
rect 1234 -109 1240 131
rect 1246 -109 1252 131
rect 1258 -109 1264 131
rect 1270 -109 1276 131
rect 1282 -109 1288 131
rect 1294 -109 1300 131
rect 1306 -109 1312 131
rect 1318 -109 1324 131
rect 1330 -109 1336 131
rect 1342 -109 1348 131
rect 1354 -109 1360 131
rect 1366 -109 1372 131
rect 1378 -109 1384 131
rect 1390 -109 1396 131
rect 1402 -109 1408 131
rect 1414 -109 1420 131
rect 1426 -109 1432 131
rect 1438 -109 1444 131
rect 1450 -109 1456 131
rect 1462 -109 1468 131
rect 1474 -109 1480 131
rect 1486 -109 1492 131
rect 1498 -109 1504 131
rect 1510 -109 1516 131
rect 1522 -109 1528 131
rect 1534 -109 1540 131
rect 1546 -109 1552 131
rect 1558 -109 1564 131
rect 1570 -109 1576 131
rect 1582 -109 1588 131
rect 1594 -109 1600 131
rect 1606 -109 1612 131
<< ndiffusion >>
rect 237 -367 238 -127
rect 242 -367 243 -127
rect 249 -367 250 -127
rect 254 -367 255 -127
rect 261 -367 262 -127
rect 266 -367 267 -127
rect 273 -367 274 -127
rect 278 -367 279 -127
rect 285 -367 286 -127
rect 290 -367 291 -127
rect 297 -367 298 -127
rect 302 -367 303 -127
rect 309 -367 310 -127
rect 314 -367 315 -127
rect 321 -367 322 -127
rect 326 -367 327 -127
rect 333 -367 334 -127
rect 338 -367 339 -127
rect 345 -367 346 -127
rect 350 -367 351 -127
rect 357 -367 358 -127
rect 362 -367 363 -127
rect 369 -367 370 -127
rect 374 -367 375 -127
rect 381 -367 382 -127
rect 386 -367 387 -127
rect 393 -367 394 -127
rect 398 -367 399 -127
rect 405 -367 406 -127
rect 410 -367 411 -127
rect 417 -367 418 -127
rect 422 -367 423 -127
rect 429 -367 430 -127
rect 434 -367 435 -127
rect 441 -367 442 -127
rect 446 -367 447 -127
rect 453 -367 454 -127
rect 458 -367 459 -127
rect 465 -367 466 -127
rect 470 -367 471 -127
rect 477 -367 478 -127
rect 482 -367 483 -127
rect 489 -367 490 -127
rect 494 -367 495 -127
rect 501 -367 502 -127
rect 506 -367 507 -127
rect 513 -367 514 -127
rect 518 -367 519 -127
rect 525 -367 526 -127
rect 530 -367 531 -127
rect 537 -367 538 -127
rect 542 -367 543 -127
rect 549 -367 550 -127
rect 554 -367 555 -127
rect 561 -367 562 -127
rect 566 -367 567 -127
rect 573 -367 574 -127
rect 578 -367 579 -127
rect 585 -367 586 -127
rect 590 -367 591 -127
rect 597 -367 598 -127
rect 602 -367 603 -127
rect 609 -367 610 -127
rect 614 -367 615 -127
rect 621 -367 622 -127
rect 626 -367 627 -127
rect 633 -367 634 -127
rect 638 -367 639 -127
rect 645 -367 646 -127
rect 650 -367 651 -127
rect 657 -367 658 -127
rect 662 -367 663 -127
rect 669 -367 670 -127
rect 674 -367 675 -127
rect 681 -367 682 -127
rect 686 -367 687 -127
rect 693 -367 694 -127
rect 698 -367 699 -127
rect 705 -367 706 -127
rect 710 -367 711 -127
rect 717 -367 718 -127
rect 722 -367 723 -127
rect 729 -367 730 -127
rect 734 -367 735 -127
rect 741 -367 742 -127
rect 746 -367 747 -127
rect 753 -367 754 -127
rect 758 -367 759 -127
rect 765 -367 766 -127
rect 770 -367 771 -127
rect 777 -367 778 -127
rect 782 -367 783 -127
rect 789 -367 790 -127
rect 794 -367 795 -127
rect 801 -367 802 -127
rect 806 -367 807 -127
rect 813 -367 814 -127
rect 818 -367 819 -127
rect 825 -367 826 -127
rect 830 -367 831 -127
rect 837 -367 838 -127
rect 842 -367 843 -127
rect 849 -367 850 -127
rect 854 -367 855 -127
rect 861 -367 862 -127
rect 866 -367 867 -127
rect 873 -367 874 -127
rect 878 -367 879 -127
rect 885 -367 886 -127
rect 890 -367 891 -127
rect 897 -367 898 -127
rect 902 -367 903 -127
rect 909 -367 910 -127
rect 914 -367 915 -127
rect 921 -367 922 -127
rect 926 -367 927 -127
rect 933 -367 934 -127
rect 938 -367 939 -127
rect 945 -367 946 -127
rect 950 -367 951 -127
rect 957 -367 958 -127
rect 962 -367 963 -127
rect 969 -367 970 -127
rect 974 -367 975 -127
rect 981 -367 982 -127
rect 986 -367 987 -127
rect 993 -367 994 -127
rect 998 -367 999 -127
rect 1005 -367 1006 -127
rect 1010 -367 1011 -127
rect 1017 -367 1018 -127
rect 1022 -367 1023 -127
rect 1029 -367 1030 -127
rect 1034 -367 1035 -127
rect 1041 -367 1042 -127
rect 1046 -367 1047 -127
rect 1053 -367 1054 -127
rect 1058 -367 1059 -127
rect 1065 -367 1066 -127
rect 1070 -367 1071 -127
rect 1077 -367 1078 -127
rect 1082 -367 1083 -127
rect 1089 -367 1090 -127
rect 1094 -367 1095 -127
rect 1101 -367 1102 -127
rect 1106 -367 1107 -127
rect 1113 -367 1114 -127
rect 1118 -367 1119 -127
rect 1125 -367 1126 -127
rect 1130 -367 1131 -127
rect 1137 -367 1138 -127
rect 1142 -367 1143 -127
rect 1149 -367 1150 -127
rect 1154 -367 1155 -127
rect 1161 -367 1162 -127
rect 1166 -367 1167 -127
rect 1173 -367 1174 -127
rect 1178 -367 1179 -127
rect 1185 -367 1186 -127
rect 1190 -367 1191 -127
rect 1197 -367 1198 -127
rect 1202 -367 1203 -127
rect 1209 -367 1210 -127
rect 1214 -367 1215 -127
rect 1221 -367 1222 -127
rect 1226 -367 1227 -127
rect 1233 -367 1234 -127
rect 1238 -367 1239 -127
rect 1245 -367 1246 -127
rect 1250 -367 1251 -127
rect 1257 -367 1258 -127
rect 1262 -367 1263 -127
rect 1269 -367 1270 -127
rect 1274 -367 1275 -127
rect 1281 -367 1282 -127
rect 1286 -367 1287 -127
rect 1293 -367 1294 -127
rect 1298 -367 1299 -127
rect 1305 -367 1306 -127
rect 1310 -367 1311 -127
rect 1317 -367 1318 -127
rect 1322 -367 1323 -127
rect 1329 -367 1330 -127
rect 1334 -367 1335 -127
rect 1341 -367 1342 -127
rect 1346 -367 1347 -127
rect 1353 -367 1354 -127
rect 1358 -367 1359 -127
rect 1365 -367 1366 -127
rect 1370 -367 1371 -127
rect 1377 -367 1378 -127
rect 1382 -367 1383 -127
rect 1389 -367 1390 -127
rect 1394 -367 1395 -127
rect 1401 -367 1402 -127
rect 1406 -367 1407 -127
rect 1413 -367 1414 -127
rect 1418 -367 1419 -127
rect 1425 -367 1426 -127
rect 1430 -367 1431 -127
rect 1437 -367 1438 -127
rect 1442 -367 1443 -127
<< pdiffusion >>
rect 237 -109 238 131
rect 242 -109 243 131
rect 249 -109 250 131
rect 254 -109 255 131
rect 261 -109 262 131
rect 266 -109 267 131
rect 273 -109 274 131
rect 278 -109 279 131
rect 285 -109 286 131
rect 290 -109 291 131
rect 297 -109 298 131
rect 302 -109 303 131
rect 309 -109 310 131
rect 314 -109 315 131
rect 321 -109 322 131
rect 326 -109 327 131
rect 333 -109 334 131
rect 338 -109 339 131
rect 345 -109 346 131
rect 350 -109 351 131
rect 357 -109 358 131
rect 362 -109 363 131
rect 369 -109 370 131
rect 374 -109 375 131
rect 381 -109 382 131
rect 386 -109 387 131
rect 393 -109 394 131
rect 398 -109 399 131
rect 405 -109 406 131
rect 410 -109 411 131
rect 417 -109 418 131
rect 422 -109 423 131
rect 429 -109 430 131
rect 434 -109 435 131
rect 441 -109 442 131
rect 446 -109 447 131
rect 453 -109 454 131
rect 458 -109 459 131
rect 465 -109 466 131
rect 470 -109 471 131
rect 477 -109 478 131
rect 482 -109 483 131
rect 489 -109 490 131
rect 494 -109 495 131
rect 501 -109 502 131
rect 506 -109 507 131
rect 513 -109 514 131
rect 518 -109 519 131
rect 525 -109 526 131
rect 530 -109 531 131
rect 537 -109 538 131
rect 542 -109 543 131
rect 549 -109 550 131
rect 554 -109 555 131
rect 561 -109 562 131
rect 566 -109 567 131
rect 573 -109 574 131
rect 578 -109 579 131
rect 585 -109 586 131
rect 590 -109 591 131
rect 597 -109 598 131
rect 602 -109 603 131
rect 609 -109 610 131
rect 614 -109 615 131
rect 621 -109 622 131
rect 626 -109 627 131
rect 633 -109 634 131
rect 638 -109 639 131
rect 645 -109 646 131
rect 650 -109 651 131
rect 657 -109 658 131
rect 662 -109 663 131
rect 669 -109 670 131
rect 674 -109 675 131
rect 681 -109 682 131
rect 686 -109 687 131
rect 693 -109 694 131
rect 698 -109 699 131
rect 705 -109 706 131
rect 710 -109 711 131
rect 717 -109 718 131
rect 722 -109 723 131
rect 729 -109 730 131
rect 734 -109 735 131
rect 741 -109 742 131
rect 746 -109 747 131
rect 753 -109 754 131
rect 758 -109 759 131
rect 765 -109 766 131
rect 770 -109 771 131
rect 777 -109 778 131
rect 782 -109 783 131
rect 789 -109 790 131
rect 794 -109 795 131
rect 801 -109 802 131
rect 806 -109 807 131
rect 813 -109 814 131
rect 818 -109 819 131
rect 825 -109 826 131
rect 830 -109 831 131
rect 837 -109 838 131
rect 842 -109 843 131
rect 1012 -109 1013 131
rect 1017 -109 1018 131
rect 1024 -109 1025 131
rect 1029 -109 1030 131
rect 1036 -109 1037 131
rect 1041 -109 1042 131
rect 1048 -109 1049 131
rect 1053 -109 1054 131
rect 1060 -109 1061 131
rect 1065 -109 1066 131
rect 1072 -109 1073 131
rect 1077 -109 1078 131
rect 1084 -109 1085 131
rect 1089 -109 1090 131
rect 1096 -109 1097 131
rect 1101 -109 1102 131
rect 1108 -109 1109 131
rect 1113 -109 1114 131
rect 1120 -109 1121 131
rect 1125 -109 1126 131
rect 1132 -109 1133 131
rect 1137 -109 1138 131
rect 1144 -109 1145 131
rect 1149 -109 1150 131
rect 1156 -109 1157 131
rect 1161 -109 1162 131
rect 1168 -109 1169 131
rect 1173 -109 1174 131
rect 1180 -109 1181 131
rect 1185 -109 1186 131
rect 1192 -109 1193 131
rect 1197 -109 1198 131
rect 1204 -109 1205 131
rect 1209 -109 1210 131
rect 1216 -109 1217 131
rect 1221 -109 1222 131
rect 1228 -109 1229 131
rect 1233 -109 1234 131
rect 1240 -109 1241 131
rect 1245 -109 1246 131
rect 1252 -109 1253 131
rect 1257 -109 1258 131
rect 1264 -109 1265 131
rect 1269 -109 1270 131
rect 1276 -109 1277 131
rect 1281 -109 1282 131
rect 1288 -109 1289 131
rect 1293 -109 1294 131
rect 1300 -109 1301 131
rect 1305 -109 1306 131
rect 1312 -109 1313 131
rect 1317 -109 1318 131
rect 1324 -109 1325 131
rect 1329 -109 1330 131
rect 1336 -109 1337 131
rect 1341 -109 1342 131
rect 1348 -109 1349 131
rect 1353 -109 1354 131
rect 1360 -109 1361 131
rect 1365 -109 1366 131
rect 1372 -109 1373 131
rect 1377 -109 1378 131
rect 1384 -109 1385 131
rect 1389 -109 1390 131
rect 1396 -109 1397 131
rect 1401 -109 1402 131
rect 1408 -109 1409 131
rect 1413 -109 1414 131
rect 1420 -109 1421 131
rect 1425 -109 1426 131
rect 1432 -109 1433 131
rect 1437 -109 1438 131
rect 1444 -109 1445 131
rect 1449 -109 1450 131
rect 1456 -109 1457 131
rect 1461 -109 1462 131
rect 1468 -109 1469 131
rect 1473 -109 1474 131
rect 1480 -109 1481 131
rect 1485 -109 1486 131
rect 1492 -109 1493 131
rect 1497 -109 1498 131
rect 1504 -109 1505 131
rect 1509 -109 1510 131
rect 1516 -109 1517 131
rect 1521 -109 1522 131
rect 1528 -109 1529 131
rect 1533 -109 1534 131
rect 1540 -109 1541 131
rect 1545 -109 1546 131
rect 1552 -109 1553 131
rect 1557 -109 1558 131
rect 1564 -109 1565 131
rect 1569 -109 1570 131
rect 1576 -109 1577 131
rect 1581 -109 1582 131
rect 1588 -109 1589 131
rect 1593 -109 1594 131
rect 1600 -109 1601 131
rect 1605 -109 1606 131
rect 1612 -109 1613 131
rect 1617 -109 1618 131
<< ndcontact >>
rect 238 -367 242 -127
rect 250 -367 254 -127
rect 262 -367 266 -127
rect 274 -367 278 -127
rect 286 -367 290 -127
rect 298 -367 302 -127
rect 310 -367 314 -127
rect 322 -367 326 -127
rect 334 -367 338 -127
rect 346 -367 350 -127
rect 358 -367 362 -127
rect 370 -367 374 -127
rect 382 -367 386 -127
rect 394 -367 398 -127
rect 406 -367 410 -127
rect 418 -367 422 -127
rect 430 -367 434 -127
rect 442 -367 446 -127
rect 454 -367 458 -127
rect 466 -367 470 -127
rect 478 -367 482 -127
rect 490 -367 494 -127
rect 502 -367 506 -127
rect 514 -367 518 -127
rect 526 -367 530 -127
rect 538 -367 542 -127
rect 550 -367 554 -127
rect 562 -367 566 -127
rect 574 -367 578 -127
rect 586 -367 590 -127
rect 598 -367 602 -127
rect 610 -367 614 -127
rect 622 -367 626 -127
rect 634 -367 638 -127
rect 646 -367 650 -127
rect 658 -367 662 -127
rect 670 -367 674 -127
rect 682 -367 686 -127
rect 694 -367 698 -127
rect 706 -367 710 -127
rect 718 -367 722 -127
rect 730 -367 734 -127
rect 742 -367 746 -127
rect 754 -367 758 -127
rect 766 -367 770 -127
rect 778 -367 782 -127
rect 790 -367 794 -127
rect 802 -367 806 -127
rect 814 -367 818 -127
rect 826 -367 830 -127
rect 838 -367 842 -127
rect 850 -367 854 -127
rect 862 -367 866 -127
rect 874 -367 878 -127
rect 886 -367 890 -127
rect 898 -367 902 -127
rect 910 -367 914 -127
rect 922 -367 926 -127
rect 934 -367 938 -127
rect 946 -367 950 -127
rect 958 -367 962 -127
rect 970 -367 974 -127
rect 982 -367 986 -127
rect 994 -367 998 -127
rect 1006 -367 1010 -127
rect 1018 -367 1022 -127
rect 1030 -367 1034 -127
rect 1042 -367 1046 -127
rect 1054 -367 1058 -127
rect 1066 -367 1070 -127
rect 1078 -367 1082 -127
rect 1090 -367 1094 -127
rect 1102 -367 1106 -127
rect 1114 -367 1118 -127
rect 1126 -367 1130 -127
rect 1138 -367 1142 -127
rect 1150 -367 1154 -127
rect 1162 -367 1166 -127
rect 1174 -367 1178 -127
rect 1186 -367 1190 -127
rect 1198 -367 1202 -127
rect 1210 -367 1214 -127
rect 1222 -367 1226 -127
rect 1234 -367 1238 -127
rect 1246 -367 1250 -127
rect 1258 -367 1262 -127
rect 1270 -367 1274 -127
rect 1282 -367 1286 -127
rect 1294 -367 1298 -127
rect 1306 -367 1310 -127
rect 1318 -367 1322 -127
rect 1330 -367 1334 -127
rect 1342 -367 1346 -127
rect 1354 -367 1358 -127
rect 1366 -367 1370 -127
rect 1378 -367 1382 -127
rect 1390 -367 1394 -127
rect 1402 -367 1406 -127
rect 1414 -367 1418 -127
rect 1426 -367 1430 -127
rect 1438 -367 1442 -127
<< pdcontact >>
rect 11 -14 15 -10
rect 103 -14 107 -10
rect 238 -109 242 131
rect 250 -109 254 131
rect 262 -109 266 131
rect 274 -109 278 131
rect 286 -109 290 131
rect 298 -109 302 131
rect 310 -109 314 131
rect 322 -109 326 131
rect 334 -109 338 131
rect 346 -109 350 131
rect 358 -109 362 131
rect 370 -109 374 131
rect 382 -109 386 131
rect 394 -109 398 131
rect 406 -109 410 131
rect 418 -109 422 131
rect 430 -109 434 131
rect 442 -109 446 131
rect 454 -109 458 131
rect 466 -109 470 131
rect 478 -109 482 131
rect 490 -109 494 131
rect 502 -109 506 131
rect 514 -109 518 131
rect 526 -109 530 131
rect 538 -109 542 131
rect 550 -109 554 131
rect 562 -109 566 131
rect 574 -109 578 131
rect 586 -109 590 131
rect 598 -109 602 131
rect 610 -109 614 131
rect 622 -109 626 131
rect 634 -109 638 131
rect 646 -109 650 131
rect 658 -109 662 131
rect 670 -109 674 131
rect 682 -109 686 131
rect 694 -109 698 131
rect 706 -109 710 131
rect 718 -109 722 131
rect 730 -109 734 131
rect 742 -109 746 131
rect 754 -109 758 131
rect 766 -109 770 131
rect 778 -109 782 131
rect 790 -109 794 131
rect 802 -109 806 131
rect 814 -109 818 131
rect 826 -109 830 131
rect 838 -109 842 131
rect 1013 -109 1017 131
rect 1025 -109 1029 131
rect 1037 -109 1041 131
rect 1049 -109 1053 131
rect 1061 -109 1065 131
rect 1073 -109 1077 131
rect 1085 -109 1089 131
rect 1097 -109 1101 131
rect 1109 -109 1113 131
rect 1121 -109 1125 131
rect 1133 -109 1137 131
rect 1145 -109 1149 131
rect 1157 -109 1161 131
rect 1169 -109 1173 131
rect 1181 -109 1185 131
rect 1193 -109 1197 131
rect 1205 -109 1209 131
rect 1217 -109 1221 131
rect 1229 -109 1233 131
rect 1241 -109 1245 131
rect 1253 -109 1257 131
rect 1265 -109 1269 131
rect 1277 -109 1281 131
rect 1289 -109 1293 131
rect 1301 -109 1305 131
rect 1313 -109 1317 131
rect 1325 -109 1329 131
rect 1337 -109 1341 131
rect 1349 -109 1353 131
rect 1361 -109 1365 131
rect 1373 -109 1377 131
rect 1385 -109 1389 131
rect 1397 -109 1401 131
rect 1409 -109 1413 131
rect 1421 -109 1425 131
rect 1433 -109 1437 131
rect 1445 -109 1449 131
rect 1457 -109 1461 131
rect 1469 -109 1473 131
rect 1481 -109 1485 131
rect 1493 -109 1497 131
rect 1505 -109 1509 131
rect 1517 -109 1521 131
rect 1529 -109 1533 131
rect 1541 -109 1545 131
rect 1553 -109 1557 131
rect 1565 -109 1569 131
rect 1577 -109 1581 131
rect 1589 -109 1593 131
rect 1601 -109 1605 131
rect 1613 -109 1617 131
<< polysilicon >>
rect 845 138 1011 219
rect 845 134 1024 138
rect 243 131 249 134
rect 255 131 261 134
rect 267 131 273 134
rect 279 131 285 134
rect 291 131 297 134
rect 303 131 309 134
rect 315 131 321 134
rect 327 131 333 134
rect 339 131 345 134
rect 351 131 357 134
rect 363 131 369 134
rect 375 131 381 134
rect 387 131 393 134
rect 399 131 405 134
rect 411 131 417 134
rect 423 131 429 134
rect 435 131 441 134
rect 447 131 453 134
rect 459 131 465 134
rect 471 131 477 134
rect 483 131 489 134
rect 495 131 501 134
rect 507 131 513 134
rect 519 131 525 134
rect 531 131 537 134
rect 543 131 549 134
rect 555 131 561 134
rect 567 131 573 134
rect 579 131 585 134
rect 591 131 597 134
rect 603 131 609 134
rect 615 131 621 134
rect 627 131 633 134
rect 639 131 645 134
rect 651 131 657 134
rect 663 131 669 134
rect 675 131 681 134
rect 687 131 693 134
rect 699 131 705 134
rect 711 131 717 134
rect 723 131 729 134
rect 735 131 741 134
rect 747 131 753 134
rect 759 131 765 134
rect 771 131 777 134
rect 783 131 789 134
rect 795 131 801 134
rect 807 131 813 134
rect 819 131 825 134
rect 831 131 837 134
rect 57 3 63 4
rect 109 3 115 4
rect 845 53 1011 134
rect 1018 131 1024 134
rect 1030 131 1036 134
rect 1042 131 1048 134
rect 1054 131 1060 134
rect 1066 131 1072 134
rect 1078 131 1084 134
rect 1090 131 1096 134
rect 1102 131 1108 134
rect 1114 131 1120 134
rect 1126 131 1132 134
rect 1138 131 1144 134
rect 1150 131 1156 134
rect 1162 131 1168 134
rect 1174 131 1180 134
rect 1186 131 1192 134
rect 1198 131 1204 134
rect 1210 131 1216 134
rect 1222 131 1228 134
rect 1234 131 1240 134
rect 1246 131 1252 134
rect 1258 131 1264 134
rect 1270 131 1276 134
rect 1282 131 1288 134
rect 1294 131 1300 134
rect 1306 131 1312 134
rect 1318 131 1324 134
rect 1330 131 1336 134
rect 1342 131 1348 134
rect 1354 131 1360 134
rect 1366 131 1372 134
rect 1378 131 1384 134
rect 1390 131 1396 134
rect 1402 131 1408 134
rect 1414 131 1420 134
rect 1426 131 1432 134
rect 1438 131 1444 134
rect 1450 131 1456 134
rect 1462 131 1468 134
rect 1474 131 1480 134
rect 1486 131 1492 134
rect 1498 131 1504 134
rect 1510 131 1516 134
rect 1522 131 1528 134
rect 1534 131 1540 134
rect 1546 131 1552 134
rect 1558 131 1564 134
rect 1570 131 1576 134
rect 1582 131 1588 134
rect 1594 131 1600 134
rect 1606 131 1612 134
rect 243 -112 249 -109
rect 255 -112 261 -109
rect 267 -112 273 -109
rect 279 -112 285 -109
rect 291 -112 297 -109
rect 303 -112 309 -109
rect 315 -112 321 -109
rect 327 -112 333 -109
rect 339 -112 345 -109
rect 351 -112 357 -109
rect 363 -112 369 -109
rect 375 -112 381 -109
rect 387 -112 393 -109
rect 399 -112 405 -109
rect 411 -112 417 -109
rect 423 -112 429 -109
rect 435 -112 441 -109
rect 447 -112 453 -109
rect 459 -112 465 -109
rect 471 -112 477 -109
rect 483 -112 489 -109
rect 495 -112 501 -109
rect 507 -112 513 -109
rect 519 -112 525 -109
rect 531 -112 537 -109
rect 543 -112 549 -109
rect 555 -112 561 -109
rect 567 -112 573 -109
rect 579 -112 585 -109
rect 591 -112 597 -109
rect 603 -112 609 -109
rect 615 -112 621 -109
rect 627 -112 633 -109
rect 639 -112 645 -109
rect 651 -112 657 -109
rect 663 -112 669 -109
rect 675 -112 681 -109
rect 687 -112 693 -109
rect 699 -112 705 -109
rect 711 -112 717 -109
rect 723 -112 729 -109
rect 735 -112 741 -109
rect 747 -112 753 -109
rect 759 -112 765 -109
rect 771 -112 777 -109
rect 783 -112 789 -109
rect 795 -112 801 -109
rect 807 -112 813 -109
rect 819 -112 825 -109
rect 831 -112 837 -109
rect 845 -112 1011 50
rect 238 -116 1011 -112
rect 1018 -112 1024 -109
rect 1030 -112 1036 -109
rect 1042 -112 1048 -109
rect 1054 -112 1060 -109
rect 1066 -112 1072 -109
rect 1078 -112 1084 -109
rect 1090 -112 1096 -109
rect 1102 -112 1108 -109
rect 1114 -112 1120 -109
rect 1126 -112 1132 -109
rect 1138 -112 1144 -109
rect 1150 -112 1156 -109
rect 1162 -112 1168 -109
rect 1174 -112 1180 -109
rect 1186 -112 1192 -109
rect 1198 -112 1204 -109
rect 1210 -112 1216 -109
rect 1222 -112 1228 -109
rect 1234 -112 1240 -109
rect 1246 -112 1252 -109
rect 1258 -112 1264 -109
rect 1270 -112 1276 -109
rect 1282 -112 1288 -109
rect 1294 -112 1300 -109
rect 1306 -112 1312 -109
rect 1318 -112 1324 -109
rect 1330 -112 1336 -109
rect 1342 -112 1348 -109
rect 1354 -112 1360 -109
rect 1366 -112 1372 -109
rect 1378 -112 1384 -109
rect 1390 -112 1396 -109
rect 1402 -112 1408 -109
rect 1414 -112 1420 -109
rect 1426 -112 1432 -109
rect 1438 -112 1444 -109
rect 1450 -112 1456 -109
rect 1462 -112 1468 -109
rect 1474 -112 1480 -109
rect 1486 -112 1492 -109
rect 1498 -112 1504 -109
rect 1510 -112 1516 -109
rect 1522 -112 1528 -109
rect 1534 -112 1540 -109
rect 1546 -112 1552 -109
rect 1558 -112 1564 -109
rect 1570 -112 1576 -109
rect 1582 -112 1588 -109
rect 1594 -112 1600 -109
rect 1606 -112 1612 -109
rect 1018 -116 1612 -112
rect 243 -127 249 -124
rect 255 -127 261 -124
rect 267 -127 273 -124
rect 279 -127 285 -124
rect 291 -127 297 -124
rect 303 -127 309 -124
rect 315 -127 321 -124
rect 327 -127 333 -124
rect 339 -127 345 -124
rect 351 -127 357 -124
rect 363 -127 369 -124
rect 375 -127 381 -124
rect 387 -127 393 -124
rect 399 -127 405 -124
rect 411 -127 417 -124
rect 423 -127 429 -124
rect 435 -127 441 -124
rect 447 -127 453 -124
rect 459 -127 465 -124
rect 471 -127 477 -124
rect 483 -127 489 -124
rect 495 -127 501 -124
rect 507 -127 513 -124
rect 519 -127 525 -124
rect 531 -127 537 -124
rect 543 -127 549 -124
rect 555 -127 561 -124
rect 567 -127 573 -124
rect 579 -127 585 -124
rect 591 -127 597 -124
rect 603 -127 609 -124
rect 615 -127 621 -124
rect 627 -127 633 -124
rect 639 -127 645 -124
rect 651 -127 657 -124
rect 663 -127 669 -124
rect 675 -127 681 -124
rect 687 -127 693 -124
rect 699 -127 705 -124
rect 711 -127 717 -124
rect 723 -127 729 -124
rect 735 -127 741 -124
rect 747 -127 753 -124
rect 759 -127 765 -124
rect 771 -127 777 -124
rect 783 -127 789 -124
rect 795 -127 801 -124
rect 807 -127 813 -124
rect 819 -127 825 -124
rect 831 -127 837 -124
rect 843 -127 849 -124
rect 855 -127 861 -124
rect 867 -127 873 -124
rect 879 -127 885 -124
rect 891 -127 897 -124
rect 903 -127 909 -124
rect 915 -127 921 -124
rect 927 -127 933 -124
rect 939 -127 945 -124
rect 951 -127 957 -124
rect 963 -127 969 -124
rect 975 -127 981 -124
rect 987 -127 993 -124
rect 999 -127 1005 -124
rect 1011 -127 1017 -124
rect 1023 -127 1029 -124
rect 1035 -127 1041 -124
rect 1047 -127 1053 -124
rect 1059 -127 1065 -124
rect 1071 -127 1077 -124
rect 1083 -127 1089 -124
rect 1095 -127 1101 -124
rect 1107 -127 1113 -124
rect 1119 -127 1125 -124
rect 1131 -127 1137 -124
rect 1143 -127 1149 -124
rect 1155 -127 1161 -124
rect 1167 -127 1173 -124
rect 1179 -127 1185 -124
rect 1191 -127 1197 -124
rect 1203 -127 1209 -124
rect 1215 -127 1221 -124
rect 1227 -127 1233 -124
rect 1239 -127 1245 -124
rect 1251 -127 1257 -124
rect 1263 -127 1269 -124
rect 1275 -127 1281 -124
rect 1287 -127 1293 -124
rect 1299 -127 1305 -124
rect 1311 -127 1317 -124
rect 1323 -127 1329 -124
rect 1335 -127 1341 -124
rect 1347 -127 1353 -124
rect 1359 -127 1365 -124
rect 1371 -127 1377 -124
rect 1383 -127 1389 -124
rect 1395 -127 1401 -124
rect 1407 -127 1413 -124
rect 1419 -127 1425 -124
rect 1431 -127 1437 -124
rect 243 -370 249 -367
rect 255 -370 261 -367
rect 267 -370 273 -367
rect 279 -370 285 -367
rect 291 -370 297 -367
rect 303 -370 309 -367
rect 315 -370 321 -367
rect 327 -370 333 -367
rect 339 -370 345 -367
rect 351 -370 357 -367
rect 363 -370 369 -367
rect 375 -370 381 -367
rect 387 -370 393 -367
rect 399 -370 405 -367
rect 411 -370 417 -367
rect 423 -370 429 -367
rect 435 -370 441 -367
rect 447 -370 453 -367
rect 459 -370 465 -367
rect 471 -370 477 -367
rect 483 -370 489 -367
rect 495 -370 501 -367
rect 507 -370 513 -367
rect 519 -370 525 -367
rect 531 -370 537 -367
rect 543 -370 549 -367
rect 555 -370 561 -367
rect 567 -370 573 -367
rect 579 -370 585 -367
rect 591 -370 597 -367
rect 603 -370 609 -367
rect 615 -370 621 -367
rect 627 -370 633 -367
rect 639 -370 645 -367
rect 651 -370 657 -367
rect 663 -370 669 -367
rect 675 -370 681 -367
rect 687 -370 693 -367
rect 699 -370 705 -367
rect 711 -370 717 -367
rect 723 -370 729 -367
rect 735 -370 741 -367
rect 747 -370 753 -367
rect 759 -370 765 -367
rect 771 -370 777 -367
rect 783 -370 789 -367
rect 795 -370 801 -367
rect 807 -370 813 -367
rect 819 -370 825 -367
rect 831 -370 837 -367
rect 237 -374 837 -370
rect 843 -370 849 -367
rect 855 -370 861 -367
rect 867 -370 873 -367
rect 879 -370 885 -367
rect 891 -370 897 -367
rect 903 -370 909 -367
rect 915 -370 921 -367
rect 927 -370 933 -367
rect 939 -370 945 -367
rect 951 -370 957 -367
rect 963 -370 969 -367
rect 975 -370 981 -367
rect 987 -370 993 -367
rect 999 -370 1005 -367
rect 1011 -370 1017 -367
rect 1023 -370 1029 -367
rect 1035 -370 1041 -367
rect 1047 -370 1053 -367
rect 1059 -370 1065 -367
rect 1071 -370 1077 -367
rect 1083 -370 1089 -367
rect 1095 -370 1101 -367
rect 1107 -370 1113 -367
rect 1119 -370 1125 -367
rect 1131 -370 1137 -367
rect 1143 -370 1149 -367
rect 1155 -370 1161 -367
rect 1167 -370 1173 -367
rect 1179 -370 1185 -367
rect 1191 -370 1197 -367
rect 1203 -370 1209 -367
rect 1215 -370 1221 -367
rect 1227 -370 1233 -367
rect 1239 -370 1245 -367
rect 1251 -370 1257 -367
rect 1263 -370 1269 -367
rect 1275 -370 1281 -367
rect 1287 -370 1293 -367
rect 1299 -370 1305 -367
rect 1311 -370 1317 -367
rect 1323 -370 1329 -367
rect 1335 -370 1341 -367
rect 1347 -370 1353 -367
rect 1359 -370 1365 -367
rect 1371 -370 1377 -367
rect 1383 -370 1389 -367
rect 1395 -370 1401 -367
rect 1407 -370 1413 -367
rect 1419 -370 1425 -367
rect 1431 -370 1437 -367
rect 843 -374 1437 -370
<< polycontact >>
rect 26 1 30 5
rect 58 -1 62 3
rect 110 -1 114 3
rect 142 1 146 5
rect 153 -9 157 -5
rect 243 -124 249 -120
rect 255 -124 261 -120
rect 267 -124 273 -120
rect 279 -124 285 -120
rect 291 -124 297 -120
rect 303 -124 309 -120
rect 315 -124 321 -120
rect 327 -124 333 -120
rect 339 -124 345 -120
rect 351 -124 357 -120
rect 363 -124 369 -120
rect 375 -124 381 -120
rect 387 -124 393 -120
rect 399 -124 405 -120
rect 411 -124 417 -120
rect 423 -124 429 -120
rect 435 -124 441 -120
rect 447 -124 453 -120
rect 459 -124 465 -120
rect 471 -124 477 -120
rect 483 -124 489 -120
rect 495 -124 501 -120
rect 507 -124 513 -120
rect 519 -124 525 -120
rect 531 -124 537 -120
rect 543 -124 549 -120
rect 555 -124 561 -120
rect 567 -124 573 -120
rect 579 -124 585 -120
rect 591 -124 597 -120
rect 603 -124 609 -120
rect 615 -124 621 -120
rect 627 -124 633 -120
rect 639 -124 645 -120
rect 651 -124 657 -120
rect 663 -124 669 -120
rect 675 -124 681 -120
rect 687 -124 693 -120
rect 699 -124 705 -120
rect 711 -124 717 -120
rect 723 -124 729 -120
rect 735 -124 741 -120
rect 747 -124 753 -120
rect 759 -124 765 -120
rect 771 -124 777 -120
rect 783 -124 789 -120
rect 795 -124 801 -120
rect 807 -124 813 -120
rect 819 -124 825 -120
rect 831 -124 837 -120
<< metal1 >>
rect 250 134 837 138
rect 250 131 254 134
rect 274 131 278 134
rect 298 131 302 134
rect 322 131 326 134
rect 346 131 350 134
rect 370 131 374 134
rect 394 131 398 134
rect 418 131 422 134
rect 442 131 446 134
rect 466 131 470 134
rect 490 131 494 134
rect 514 131 518 134
rect 538 131 542 134
rect 562 131 566 134
rect 586 131 590 134
rect 610 131 614 134
rect 634 131 638 134
rect 658 131 662 134
rect 682 131 686 134
rect 706 131 710 134
rect 730 131 734 134
rect 754 131 758 134
rect 778 131 782 134
rect 802 131 806 134
rect 826 131 830 134
rect 26 -1 30 1
rect 11 -5 30 -1
rect 58 -5 62 -1
rect 103 -5 114 -1
rect 142 0 146 1
rect 142 -4 157 0
rect 153 -5 157 -4
rect 11 -10 15 -5
rect 103 -10 107 -5
rect 1025 134 1605 138
rect 1025 131 1029 134
rect 1049 131 1053 134
rect 1073 131 1077 134
rect 1097 131 1101 134
rect 1121 131 1125 134
rect 1145 131 1149 134
rect 1169 131 1173 134
rect 1193 131 1197 134
rect 1217 131 1221 134
rect 1241 131 1245 134
rect 1265 131 1269 134
rect 1289 131 1293 134
rect 1313 131 1317 134
rect 1337 131 1341 134
rect 1361 131 1365 134
rect 1385 131 1389 134
rect 1409 131 1413 134
rect 1433 131 1437 134
rect 1457 131 1461 134
rect 1481 131 1485 134
rect 1505 131 1509 134
rect 1529 131 1533 134
rect 1553 131 1557 134
rect 1577 131 1581 134
rect 1601 131 1605 134
rect 238 -112 242 -109
rect 262 -112 266 -109
rect 286 -112 290 -109
rect 310 -112 314 -109
rect 334 -112 338 -109
rect 358 -112 362 -109
rect 382 -112 386 -109
rect 406 -112 410 -109
rect 430 -112 434 -109
rect 454 -112 458 -109
rect 478 -112 482 -109
rect 502 -112 506 -109
rect 526 -112 530 -109
rect 550 -112 554 -109
rect 574 -112 578 -109
rect 598 -112 602 -109
rect 622 -112 626 -109
rect 646 -112 650 -109
rect 670 -112 674 -109
rect 694 -112 698 -109
rect 718 -112 722 -109
rect 742 -112 746 -109
rect 766 -112 770 -109
rect 790 -112 794 -109
rect 814 -112 818 -109
rect 838 -112 842 -109
rect 852 -112 856 -107
rect 238 -116 856 -112
rect 1000 -112 1004 60
rect 1013 -112 1017 -109
rect 1037 -112 1041 -109
rect 1061 -112 1065 -109
rect 1085 -112 1089 -109
rect 1109 -112 1113 -109
rect 1133 -112 1137 -109
rect 1157 -112 1161 -109
rect 1181 -112 1185 -109
rect 1205 -112 1209 -109
rect 1229 -112 1233 -109
rect 1253 -112 1257 -109
rect 1277 -112 1281 -109
rect 1301 -112 1305 -109
rect 1325 -112 1329 -109
rect 1349 -112 1353 -109
rect 1373 -112 1377 -109
rect 1397 -112 1401 -109
rect 1421 -112 1425 -109
rect 1445 -112 1449 -109
rect 1469 -112 1473 -109
rect 1493 -112 1497 -109
rect 1517 -112 1521 -109
rect 1541 -112 1545 -109
rect 1565 -112 1569 -109
rect 1589 -112 1593 -109
rect 1613 -112 1617 -109
rect 1000 -116 1617 -112
rect 243 -120 837 -116
rect 1000 -120 1430 -116
rect 249 -124 255 -120
rect 261 -124 267 -120
rect 273 -124 279 -120
rect 285 -124 291 -120
rect 297 -124 303 -120
rect 309 -124 315 -120
rect 321 -124 327 -120
rect 333 -124 339 -120
rect 345 -124 351 -120
rect 357 -124 363 -120
rect 369 -124 375 -120
rect 381 -124 387 -120
rect 393 -124 399 -120
rect 405 -124 411 -120
rect 417 -124 423 -120
rect 429 -124 435 -120
rect 441 -124 447 -120
rect 453 -124 459 -120
rect 465 -124 471 -120
rect 477 -124 483 -120
rect 489 -124 495 -120
rect 501 -124 507 -120
rect 513 -124 519 -120
rect 525 -124 531 -120
rect 537 -124 543 -120
rect 549 -124 555 -120
rect 561 -124 567 -120
rect 573 -124 579 -120
rect 585 -124 591 -120
rect 597 -124 603 -120
rect 609 -124 615 -120
rect 621 -124 627 -120
rect 633 -124 639 -120
rect 645 -124 651 -120
rect 657 -124 663 -120
rect 669 -124 675 -120
rect 681 -124 687 -120
rect 693 -124 699 -120
rect 705 -124 711 -120
rect 717 -124 723 -120
rect 729 -124 735 -120
rect 741 -124 747 -120
rect 753 -124 759 -120
rect 765 -124 771 -120
rect 777 -124 783 -120
rect 789 -124 795 -120
rect 801 -124 807 -120
rect 813 -124 819 -120
rect 825 -124 831 -120
rect 850 -124 1430 -120
rect 250 -127 254 -124
rect 274 -127 278 -124
rect 298 -127 302 -124
rect 322 -127 326 -124
rect 346 -127 350 -124
rect 370 -127 374 -124
rect 394 -127 398 -124
rect 418 -127 422 -124
rect 442 -127 446 -124
rect 466 -127 470 -124
rect 490 -127 494 -124
rect 514 -127 518 -124
rect 538 -127 542 -124
rect 562 -127 566 -124
rect 586 -127 590 -124
rect 610 -127 614 -124
rect 634 -127 638 -124
rect 658 -127 662 -124
rect 682 -127 686 -124
rect 706 -127 710 -124
rect 730 -127 734 -124
rect 754 -127 758 -124
rect 778 -127 782 -124
rect 802 -127 806 -124
rect 826 -127 830 -124
rect 850 -127 854 -124
rect 874 -127 878 -124
rect 898 -127 902 -124
rect 922 -127 926 -124
rect 946 -127 950 -124
rect 970 -127 974 -124
rect 994 -127 998 -124
rect 1018 -127 1022 -124
rect 1042 -127 1046 -124
rect 1066 -127 1070 -124
rect 1090 -127 1094 -124
rect 1114 -127 1118 -124
rect 1138 -127 1142 -124
rect 1162 -127 1166 -124
rect 1186 -127 1190 -124
rect 1210 -127 1214 -124
rect 1234 -127 1238 -124
rect 1258 -127 1262 -124
rect 1282 -127 1286 -124
rect 1306 -127 1310 -124
rect 1330 -127 1334 -124
rect 1354 -127 1358 -124
rect 1378 -127 1382 -124
rect 1402 -127 1406 -124
rect 1426 -127 1430 -124
rect 238 -370 242 -367
rect 262 -370 266 -367
rect 286 -370 290 -367
rect 310 -370 314 -367
rect 334 -370 338 -367
rect 358 -370 362 -367
rect 382 -370 386 -367
rect 406 -370 410 -367
rect 430 -370 434 -367
rect 454 -370 458 -367
rect 478 -370 482 -367
rect 502 -370 506 -367
rect 526 -370 530 -367
rect 550 -370 554 -367
rect 574 -370 578 -367
rect 598 -370 602 -367
rect 622 -370 626 -367
rect 646 -370 650 -367
rect 670 -370 674 -367
rect 694 -370 698 -367
rect 718 -370 722 -367
rect 742 -370 746 -367
rect 766 -370 770 -367
rect 790 -370 794 -367
rect 814 -370 818 -367
rect 838 -370 842 -367
rect 862 -370 866 -367
rect 886 -370 890 -367
rect 910 -370 914 -367
rect 934 -370 938 -367
rect 958 -370 962 -367
rect 982 -370 986 -367
rect 1006 -370 1010 -367
rect 1030 -370 1034 -367
rect 1054 -370 1058 -367
rect 1078 -370 1082 -367
rect 1102 -370 1106 -367
rect 1126 -370 1130 -367
rect 1150 -370 1154 -367
rect 1174 -370 1178 -367
rect 1198 -370 1202 -367
rect 1222 -370 1226 -367
rect 1246 -370 1250 -367
rect 1270 -370 1274 -367
rect 1294 -370 1298 -367
rect 1318 -370 1322 -367
rect 1342 -370 1346 -367
rect 1366 -370 1370 -367
rect 1390 -370 1394 -367
rect 1414 -370 1418 -367
rect 1438 -370 1442 -367
rect 237 -374 1442 -370
use amp  amp_0
timestamp 1418768421
transform 1 0 95 0 1 135
box -95 -135 77 126
use bias  bias_0
timestamp 1418768461
transform 1 0 -11 0 1 -106
box 13 -282 183 102
<< labels >>
rlabel metal1 838 -374 842 -370 1 Gnd
<< end >>
