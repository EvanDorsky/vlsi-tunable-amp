magic
tech scmos
timestamp 1417991047
<< ntransistor >>
rect -5 -138 -1 -136
rect 6 -138 10 -136
rect 0 -145 4 -143
<< ptransistor >>
rect -8 -88 -5 -86
rect 1 -88 4 -86
rect -5 -108 -1 -106
rect 6 -108 10 -106
<< ndiffusion >>
rect -5 -136 -1 -135
rect 6 -136 10 -135
rect -5 -139 -1 -138
rect 6 -139 10 -138
rect -5 -142 10 -139
rect 0 -143 4 -142
rect 0 -146 4 -145
rect -1 -149 6 -146
<< pdiffusion >>
rect -8 -86 -5 -85
rect 1 -86 4 -85
rect -8 -89 -5 -88
rect 1 -89 4 -88
rect -5 -106 -1 -105
rect 6 -106 10 -105
rect -5 -109 -1 -108
rect 6 -109 10 -108
<< ndcontact >>
rect -5 -135 -1 -131
rect 6 -135 10 -131
rect -5 -150 -1 -146
rect 6 -150 10 -146
<< pdcontact >>
rect -8 -85 -4 -81
rect 0 -85 4 -81
rect -8 -93 -4 -89
rect 0 -93 4 -89
rect -5 -105 -1 -101
rect 6 -105 10 -101
rect -5 -113 -1 -109
rect 6 -113 10 -109
<< polysilicon >>
rect -11 -88 -8 -86
rect -5 -88 1 -86
rect 4 -88 16 -86
rect -8 -108 -5 -106
rect -1 -108 1 -106
rect 4 -108 6 -106
rect 10 -108 13 -106
rect -8 -126 -6 -108
rect 11 -116 13 -108
rect 3 -118 13 -116
rect -8 -128 2 -126
rect -8 -136 -6 -128
rect 11 -136 13 -118
rect -8 -138 -5 -136
rect -1 -138 1 -136
rect 4 -138 6 -136
rect 10 -138 13 -136
rect -11 -145 0 -143
rect 4 -145 16 -143
<< polycontact >>
rect -1 -119 3 -115
rect 2 -129 6 -125
<< metal1 >>
rect -11 -77 2 -74
rect -1 -81 2 -77
rect 13 -77 16 -74
rect -11 -84 -8 -81
rect -1 -85 0 -81
rect 13 -84 16 -81
rect -8 -94 -4 -93
rect 0 -94 4 -93
rect -11 -105 -5 -101
rect -1 -105 6 -101
rect 10 -105 16 -101
rect -5 -120 -1 -113
rect -5 -131 -1 -124
rect 6 -120 10 -113
rect 6 -131 10 -124
rect -11 -146 16 -145
rect -11 -149 -5 -146
rect -1 -149 6 -146
rect 10 -149 16 -146
<< m2contact >>
rect 9 -78 13 -74
rect 9 -85 13 -81
rect -8 -98 -4 -94
rect 0 -98 4 -94
rect -5 -124 -1 -120
rect 6 -124 10 -120
<< metal2 >>
rect -8 -77 9 -74
rect -8 -94 -5 -77
rect -1 -84 9 -81
rect -1 -94 2 -84
rect -1 -98 0 -94
rect -8 -124 -5 -98
rect -1 -114 2 -98
rect -1 -117 10 -114
rect 6 -120 10 -117
<< labels >>
rlabel metal1 -11 -77 -10 -74 3 Dbar
rlabel metal1 -11 -84 -10 -81 3 Dbar
rlabel metal1 15 -149 16 -145 8 Gnd
rlabel metal1 15 -84 16 -81 7 Qbar
rlabel polysilicon 15 -88 16 -86 7 Clk
rlabel metal1 15 -105 16 -101 7 Vdd
rlabel polysilicon -11 -145 -10 -143 3 Clk
rlabel metal1 15 -77 16 -74 6 Q
<< end >>
