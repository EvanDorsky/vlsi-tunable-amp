magic
tech scmos
magscale 1 3
timestamp 1419057840
<< metal1 >>
rect 3290 7350 3320 7370
rect 3280 7340 3320 7350
rect 3400 7340 3410 7350
rect 3280 7330 3310 7340
rect 3350 7330 3360 7340
rect 3120 7320 3130 7330
rect 3110 7310 3130 7320
rect 3420 7310 3440 7320
rect 2820 7300 2830 7310
rect 2980 7300 3000 7310
rect 3100 7300 3130 7310
rect 3390 7300 3450 7310
rect 3460 7300 3480 7310
rect 3520 7300 3540 7310
rect 2970 7290 3000 7300
rect 3380 7290 3440 7300
rect 3460 7290 3490 7300
rect 3500 7290 3550 7300
rect 2590 7280 2620 7290
rect 2810 7280 2820 7290
rect 2950 7280 2990 7290
rect 3370 7280 3430 7290
rect 2560 7270 2570 7280
rect 2590 7260 2610 7280
rect 2960 7270 2980 7280
rect 3360 7270 3430 7280
rect 3460 7280 3580 7290
rect 3640 7280 3650 7290
rect 3460 7270 3620 7280
rect 2960 7260 2970 7270
rect 3070 7260 3110 7270
rect 3150 7260 3190 7270
rect 3340 7260 3400 7270
rect 2510 7230 2520 7250
rect 2570 7220 2610 7260
rect 2910 7250 2930 7260
rect 3060 7250 3110 7260
rect 3140 7250 3190 7260
rect 3330 7250 3380 7260
rect 3420 7250 3650 7270
rect 2900 7240 2930 7250
rect 3000 7240 3010 7250
rect 3040 7240 3090 7250
rect 2890 7230 2920 7240
rect 3030 7239 3090 7240
rect 3130 7240 3180 7250
rect 3310 7240 3350 7250
rect 3400 7240 3660 7250
rect 3030 7230 3081 7239
rect 3130 7230 3160 7240
rect 3300 7230 3340 7240
rect 3390 7230 3660 7240
rect 2870 7220 2900 7230
rect 3000 7220 3060 7230
rect 3090 7220 3100 7230
rect 3120 7220 3150 7230
rect 3290 7220 3320 7230
rect 3380 7220 3550 7230
rect 3570 7220 3590 7230
rect 3600 7220 3670 7230
rect 3780 7220 3810 7230
rect 2570 7200 2600 7220
rect 2560 7180 2600 7200
rect 2800 7200 2820 7220
rect 2870 7210 2880 7220
rect 2940 7210 2960 7220
rect 2990 7210 3050 7220
rect 3090 7210 3150 7220
rect 3280 7210 3310 7220
rect 3360 7210 3450 7220
rect 3470 7210 3490 7220
rect 3600 7210 3620 7220
rect 3630 7210 3690 7220
rect 3740 7210 3810 7220
rect 2850 7200 2860 7210
rect 2930 7200 3040 7210
rect 3080 7200 3140 7210
rect 3280 7200 3300 7210
rect 3350 7200 3420 7210
rect 3610 7200 3620 7210
rect 3640 7200 3650 7210
rect 3710 7200 3810 7210
rect 2800 7190 2810 7200
rect 2840 7190 2860 7200
rect 2910 7190 3040 7200
rect 3050 7190 3130 7200
rect 3330 7190 3400 7200
rect 3570 7190 3580 7200
rect 3700 7190 3840 7200
rect 2770 7180 2810 7190
rect 2830 7180 2850 7190
rect 2550 7170 2590 7180
rect 2760 7170 2850 7180
rect 2900 7180 3080 7190
rect 3320 7180 3360 7190
rect 3470 7180 3490 7190
rect 3560 7180 3590 7190
rect 2900 7170 3070 7180
rect 3130 7170 3150 7180
rect 3210 7170 3230 7180
rect 3300 7170 3340 7180
rect 3460 7170 3480 7180
rect 3550 7170 3590 7180
rect 2550 7160 2570 7170
rect 2750 7160 2840 7170
rect 2470 7150 2480 7160
rect 2540 7140 2570 7160
rect 2740 7150 2840 7160
rect 2890 7160 3070 7170
rect 3110 7160 3120 7170
rect 3200 7160 3220 7170
rect 3290 7160 3320 7170
rect 3440 7160 3480 7170
rect 3510 7160 3540 7170
rect 3570 7160 3580 7170
rect 3610 7160 3630 7190
rect 3700 7180 3720 7190
rect 3730 7188 3750 7190
rect 3690 7179 3720 7180
rect 3741 7180 3750 7188
rect 3760 7180 3780 7190
rect 3741 7179 3780 7180
rect 3690 7170 3730 7179
rect 3740 7170 3780 7179
rect 3800 7179 3850 7190
rect 3800 7170 3837 7179
rect 3670 7160 3790 7170
rect 3810 7160 3837 7170
rect 2890 7158 3060 7160
rect 2890 7150 3048 7158
rect 3080 7150 3120 7160
rect 3180 7150 3210 7160
rect 3280 7150 3310 7160
rect 3440 7150 3530 7160
rect 3670 7150 3800 7160
rect 3870 7158 3880 7160
rect 3850 7150 3880 7158
rect 2710 7140 2830 7150
rect 2890 7140 3030 7150
rect 3069 7149 3130 7150
rect 3060 7140 3130 7149
rect 3170 7140 3210 7150
rect 3270 7140 3290 7150
rect 3400 7140 3410 7150
rect 3420 7140 3480 7150
rect 3490 7140 3500 7150
rect 3560 7140 3590 7150
rect 3660 7140 3810 7150
rect 3840 7140 3920 7150
rect 2360 7130 2370 7140
rect 2540 7130 2560 7140
rect 2700 7130 2820 7140
rect 2870 7130 3030 7140
rect 2330 7120 2380 7130
rect 2310 7110 2380 7120
rect 2290 7090 2380 7110
rect 2530 7100 2550 7130
rect 2700 7120 2810 7130
rect 2850 7120 3020 7130
rect 3050 7120 3110 7140
rect 3160 7130 3201 7140
rect 3150 7120 3201 7130
rect 3240 7120 3250 7140
rect 3390 7130 3470 7140
rect 3550 7130 3600 7140
rect 3660 7130 3830 7140
rect 3850 7130 3910 7140
rect 3970 7130 3990 7140
rect 3330 7120 3360 7130
rect 3380 7120 3450 7130
rect 3520 7120 3530 7130
rect 3540 7120 3600 7130
rect 2700 7100 2800 7120
rect 2840 7110 3018 7120
rect 3040 7110 3070 7120
rect 3080 7110 3110 7120
rect 3130 7110 3201 7120
rect 3210 7119 3222 7120
rect 3210 7110 3230 7119
rect 3280 7110 3290 7120
rect 3330 7110 3350 7120
rect 3370 7110 3410 7120
rect 3520 7110 3590 7120
rect 2830 7100 3018 7110
rect 3030 7100 3060 7110
rect 2520 7090 2550 7100
rect 2690 7090 2790 7100
rect 2820 7090 3070 7100
rect 3080 7090 3170 7110
rect 3190 7100 3230 7110
rect 3320 7100 3340 7110
rect 3370 7100 3400 7110
rect 3510 7100 3590 7110
rect 3650 7110 3690 7130
rect 3710 7120 3840 7130
rect 3850 7120 3900 7130
rect 3710 7110 3880 7120
rect 3960 7110 3981 7130
rect 3650 7100 3740 7110
rect 3760 7100 3870 7110
rect 3920 7100 3950 7110
rect 3970 7100 3980 7110
rect 3990 7100 4010 7110
rect 4050 7100 4060 7110
rect 3200 7092 3230 7100
rect 3200 7090 3228 7092
rect 2280 7080 2370 7090
rect 2400 7080 2410 7090
rect 2290 7070 2380 7080
rect 2400 7070 2420 7080
rect 2520 7070 2540 7090
rect 2650 7080 2800 7090
rect 2810 7080 3160 7090
rect 3190 7080 3220 7090
rect 3300 7080 3330 7100
rect 3490 7090 3590 7100
rect 3640 7090 3720 7100
rect 3760 7090 3880 7100
rect 3890 7090 3960 7100
rect 3470 7089 3590 7090
rect 3470 7080 3579 7089
rect 3760 7080 3950 7090
rect 2640 7070 3160 7080
rect 3189 7071 3220 7080
rect 3210 7070 3220 7071
rect 3290 7070 3320 7080
rect 3450 7070 3480 7080
rect 3490 7070 3560 7080
rect 2290 7050 2370 7070
rect 2260 7040 2370 7050
rect 2390 7050 2410 7070
rect 2510 7060 2540 7070
rect 2570 7060 2580 7070
rect 2510 7050 2530 7060
rect 2390 7040 2420 7050
rect 2240 7010 2360 7040
rect 2380 7020 2420 7040
rect 2470 7020 2480 7030
rect 2370 7010 2420 7020
rect 2460 7011 2480 7020
rect 2500 7010 2530 7050
rect 2560 7030 2580 7060
rect 2250 6990 2420 7010
rect 2490 6999 2530 7010
rect 2550 7000 2580 7030
rect 2640 7060 3150 7070
rect 2640 7030 2770 7060
rect 2790 7050 3150 7060
rect 3210 7068 3228 7070
rect 3210 7059 3240 7068
rect 3290 7060 3310 7070
rect 3400 7060 3470 7070
rect 3200 7050 3240 7059
rect 3280 7050 3300 7060
rect 3390 7050 3430 7060
rect 3450 7050 3460 7060
rect 3500 7050 3560 7070
rect 3590 7070 3600 7080
rect 3610 7070 3640 7080
rect 3760 7070 3780 7080
rect 3590 7060 3620 7070
rect 3680 7060 3690 7070
rect 3770 7060 3780 7070
rect 3580 7050 3610 7060
rect 3670 7050 3700 7060
rect 3760 7050 3780 7060
rect 3801 7070 3810 7080
rect 3820 7070 3870 7080
rect 3801 7060 3850 7070
rect 3990 7060 4040 7070
rect 3801 7050 3810 7060
rect 3970 7050 4080 7060
rect 2790 7040 3080 7050
rect 3090 7041 3140 7050
rect 3090 7040 3153 7041
rect 3170 7040 3180 7050
rect 3200 7040 3230 7050
rect 2780 7030 3210 7040
rect 3320 7030 3330 7050
rect 3390 7040 3420 7050
rect 3490 7040 3550 7050
rect 2640 7010 3210 7030
rect 3260 7020 3270 7030
rect 3300 7020 3330 7030
rect 3480 7030 3540 7040
rect 3570 7030 3600 7050
rect 3660 7040 3690 7050
rect 3750 7040 3780 7050
rect 3950 7040 4090 7050
rect 3660 7030 3680 7040
rect 3750 7030 3760 7040
rect 3920 7030 4100 7040
rect 3480 7020 3530 7030
rect 3570 7020 3590 7030
rect 3650 7020 3670 7030
rect 3720 7020 3730 7030
rect 3880 7020 4110 7030
rect 3290 7010 3320 7020
rect 3470 7010 3530 7020
rect 3560 7010 3590 7020
rect 3880 7010 4010 7020
rect 4030 7010 4140 7020
rect 2630 7000 3210 7010
rect 3250 7000 3260 7010
rect 2480 6990 2530 6999
rect 2240 6980 2430 6990
rect 2460 6980 2530 6990
rect 2540 6980 2580 7000
rect 2620 6990 3180 7000
rect 3189 6999 3210 7000
rect 3200 6990 3210 6999
rect 3240 6990 3260 7000
rect 3280 7000 3320 7010
rect 3280 6990 3300 7000
rect 3460 6990 3520 7010
rect 3560 6990 3580 7010
rect 3870 7000 3930 7010
rect 3860 6993 3920 7000
rect 3948 6999 4000 7010
rect 4030 7000 4150 7010
rect 3849 6990 3920 6993
rect 3950 6990 4000 6999
rect 4020 6990 4160 7000
rect 2610 6980 3210 6990
rect 3230 6980 3290 6990
rect 3450 6980 3510 6990
rect 3849 6980 3890 6990
rect 3950 6980 3990 6990
rect 4020 6980 4170 6990
rect 2250 6910 2430 6980
rect 2450 6960 2470 6980
rect 2480 6950 2520 6980
rect 2540 6970 3180 6980
rect 2540 6960 3160 6970
rect 3170 6960 3180 6970
rect 2470 6940 2520 6950
rect 2530 6950 3180 6960
rect 3200 6960 3310 6980
rect 3450 6970 3500 6980
rect 3849 6978 3873 6980
rect 3849 6970 3860 6978
rect 3950 6975 3980 6980
rect 3480 6960 3490 6970
rect 3560 6960 3570 6970
rect 3840 6963 3860 6970
rect 3200 6950 3300 6960
rect 3470 6950 3490 6960
rect 3550 6950 3570 6960
rect 3825 6960 3860 6963
rect 3939 6960 3980 6975
rect 4020 6970 4180 6980
rect 4010 6960 4170 6970
rect 3825 6950 3850 6960
rect 3920 6950 3950 6960
rect 3960 6950 3970 6960
rect 4000 6950 4120 6960
rect 4140 6950 4160 6960
rect 2530 6940 3270 6950
rect 3460 6940 3480 6950
rect 3540 6940 3560 6950
rect 3820 6948 3849 6950
rect 3820 6940 3840 6948
rect 3910 6940 3950 6950
rect 4000 6940 4110 6950
rect 2470 6920 3250 6940
rect 3370 6920 3380 6930
rect 3440 6920 3470 6940
rect 3540 6930 3550 6940
rect 3810 6930 3830 6940
rect 3910 6930 3930 6940
rect 3980 6930 4140 6940
rect 3810 6920 3820 6930
rect 3890 6920 3920 6930
rect 3980 6920 4000 6930
rect 4030 6920 4080 6930
rect 4100 6920 4130 6930
rect 4230 6920 4260 6930
rect 2470 6910 3240 6920
rect 3330 6910 3340 6920
rect 3360 6910 3380 6920
rect 3430 6910 3460 6920
rect 3870 6910 3900 6920
rect 2230 6890 2440 6910
rect 2470 6890 3230 6910
rect 3270 6900 3280 6910
rect 3320 6909 3340 6910
rect 3350 6909 3370 6910
rect 3320 6900 3370 6909
rect 3430 6900 3450 6910
rect 3860 6900 3900 6910
rect 4040 6910 4080 6920
rect 4110 6910 4130 6920
rect 4210 6910 4260 6920
rect 4040 6900 4070 6910
rect 4200 6900 4250 6910
rect 3250 6890 3280 6900
rect 2240 6880 2440 6890
rect 2250 6860 2440 6880
rect 2240 6850 2440 6860
rect 2230 6840 2440 6850
rect 2460 6870 3220 6890
rect 3240 6880 3280 6890
rect 3327 6885 3360 6900
rect 3850 6890 3900 6900
rect 3940 6890 3960 6900
rect 3990 6890 4050 6900
rect 4190 6890 4230 6900
rect 3330 6880 3360 6885
rect 3530 6880 3550 6890
rect 3780 6880 3810 6890
rect 3840 6880 3891 6890
rect 3230 6870 3270 6880
rect 3330 6870 3350 6880
rect 3420 6870 3460 6880
rect 3510 6870 3550 6880
rect 3770 6870 3800 6880
rect 3830 6879 3891 6880
rect 3930 6880 3960 6890
rect 3980 6880 4040 6890
rect 4170 6880 4210 6890
rect 3830 6870 3860 6879
rect 2460 6860 2520 6870
rect 2530 6860 3270 6870
rect 3320 6860 3350 6870
rect 3400 6860 3460 6870
rect 3490 6860 3540 6870
rect 3760 6860 3790 6870
rect 3820 6860 3850 6870
rect 3880 6860 3890 6879
rect 3930 6870 4040 6880
rect 4150 6870 4200 6880
rect 3930 6860 3990 6870
rect 4020 6860 4040 6870
rect 4140 6860 4180 6870
rect 2460 6850 3260 6860
rect 3310 6850 3350 6860
rect 3390 6850 3460 6860
rect 3470 6850 3530 6860
rect 3690 6850 3710 6860
rect 2460 6840 3250 6850
rect 2220 6830 2450 6840
rect 2230 6810 2450 6830
rect 2220 6800 2450 6810
rect 2210 6765 2450 6800
rect 2460 6830 3100 6840
rect 3120 6830 3250 6840
rect 3300 6830 3340 6850
rect 3380 6840 3520 6850
rect 3540 6840 3560 6850
rect 3370 6830 3510 6840
rect 3540 6830 3550 6840
rect 3600 6830 3620 6850
rect 3670 6840 3710 6850
rect 3750 6849 3770 6860
rect 3800 6850 3830 6860
rect 3910 6850 3980 6860
rect 3750 6840 3780 6849
rect 3790 6840 3820 6850
rect 3880 6840 3980 6850
rect 4030 6850 4050 6860
rect 4130 6850 4170 6860
rect 4350 6850 4360 6860
rect 3990 6840 4011 6843
rect 4030 6840 4040 6850
rect 4100 6840 4150 6850
rect 4350 6840 4370 6850
rect 3670 6830 3740 6840
rect 3770 6830 3810 6840
rect 3870 6830 4011 6840
rect 4020 6830 4040 6840
rect 4090 6830 4130 6840
rect 4300 6830 4320 6840
rect 4360 6830 4370 6840
rect 2460 6810 3080 6830
rect 3110 6820 3260 6830
rect 3280 6820 3290 6830
rect 2460 6800 3070 6810
rect 3110 6800 3250 6820
rect 3270 6810 3290 6820
rect 3300 6820 3330 6830
rect 3360 6820 3410 6830
rect 3420 6820 3510 6830
rect 3530 6820 3560 6830
rect 3580 6820 3740 6830
rect 3760 6820 3810 6830
rect 3880 6820 4040 6830
rect 4070 6820 4130 6830
rect 4290 6820 4310 6830
rect 3300 6810 3320 6820
rect 3350 6810 3550 6820
rect 3270 6800 3320 6810
rect 3340 6800 3490 6810
rect 3500 6800 3550 6810
rect 3570 6819 3732 6820
rect 3570 6810 3720 6819
rect 3750 6810 3810 6820
rect 3870 6810 4050 6820
rect 4060 6810 4140 6820
rect 4200 6810 4230 6820
rect 4290 6810 4300 6820
rect 3570 6807 3710 6810
rect 3570 6800 3708 6807
rect 3740 6800 4230 6810
rect 2460 6790 3080 6800
rect 3100 6790 3240 6800
rect 3260 6790 3310 6800
rect 2460 6780 3070 6790
rect 3100 6780 3210 6790
rect 3220 6780 3240 6790
rect 2460 6770 3060 6780
rect 3120 6770 3200 6780
rect 3250 6770 3310 6790
rect 3330 6790 3470 6800
rect 3500 6790 3700 6800
rect 3730 6790 3770 6800
rect 3330 6780 3360 6790
rect 3330 6770 3340 6780
rect 3370 6770 3460 6790
rect 3490 6780 3700 6790
rect 3710 6780 3770 6790
rect 3790 6790 4100 6800
rect 4110 6790 4210 6800
rect 4360 6790 4410 6800
rect 3790 6780 4190 6790
rect 4240 6780 4260 6790
rect 4360 6780 4400 6790
rect 3470 6770 4190 6780
rect 4230 6770 4260 6780
rect 4310 6770 4330 6780
rect 2210 6750 2260 6765
rect 2270 6760 2450 6765
rect 2470 6760 3050 6770
rect 2280 6750 2440 6760
rect 2470 6750 3040 6760
rect 3120 6750 3190 6770
rect 3240 6760 3310 6770
rect 3370 6760 3410 6770
rect 3450 6760 4260 6770
rect 4290 6760 4330 6770
rect 4410 6760 4440 6770
rect 3240 6750 3300 6760
rect 3370 6750 3400 6760
rect 3440 6750 4320 6760
rect 4400 6750 4440 6760
rect 2200 6740 2440 6750
rect 2460 6740 3030 6750
rect 3130 6740 3180 6750
rect 2200 6730 2840 6740
rect 2870 6730 2880 6740
rect 2970 6730 3020 6740
rect 3130 6730 3150 6740
rect 3240 6735 3280 6750
rect 3360 6740 3380 6750
rect 3420 6740 4180 6750
rect 4190 6740 4320 6750
rect 3250 6730 3280 6735
rect 3420 6730 4330 6740
rect 4370 6730 4380 6740
rect 2200 6710 2260 6730
rect 2270 6720 2820 6730
rect 3250 6720 3270 6730
rect 3420 6720 3560 6730
rect 2270 6710 2800 6720
rect 3400 6710 3450 6720
rect 3470 6710 3560 6720
rect 3570 6720 4350 6730
rect 3570 6710 4340 6720
rect 2230 6700 2740 6710
rect 2760 6700 2790 6710
rect 3400 6700 3440 6710
rect 3470 6700 3600 6710
rect 3610 6700 3650 6710
rect 3670 6700 4260 6710
rect 2240 6690 2730 6700
rect 3210 6690 3220 6700
rect 3400 6690 3410 6700
rect 3470 6690 3520 6700
rect 3550 6690 3600 6700
rect 3620 6690 3640 6700
rect 3670 6690 3800 6700
rect 2240 6680 2690 6690
rect 2700 6680 2710 6690
rect 3470 6681 3490 6690
rect 3471 6680 3490 6681
rect 3560 6680 3600 6690
rect 3680 6680 3690 6690
rect 3730 6680 3800 6690
rect 3810 6690 4260 6700
rect 4280 6700 4320 6710
rect 4280 6690 4310 6700
rect 4390 6690 4410 6700
rect 3810 6680 4310 6690
rect 2240 6670 2660 6680
rect 3471 6670 3480 6680
rect 3560 6670 3570 6680
rect 3580 6670 3590 6680
rect 3730 6670 4323 6680
rect 4360 6670 4370 6680
rect 2240 6660 2640 6670
rect 3740 6660 3850 6670
rect 3870 6660 4320 6670
rect 4350 6669 4380 6670
rect 4340 6660 4380 6669
rect 2240 6650 2610 6660
rect 3730 6650 4420 6660
rect 2240 6640 2590 6650
rect 3730 6640 4450 6650
rect 2200 6620 2210 6640
rect 2240 6630 2580 6640
rect 3720 6630 4460 6640
rect 2230 6620 2560 6630
rect 3710 6620 3780 6630
rect 3820 6620 3930 6630
rect 3970 6620 4330 6630
rect 4360 6620 4380 6630
rect 4440 6620 4461 6630
rect 2220 6610 2550 6620
rect 3720 6610 3730 6620
rect 3820 6610 3900 6620
rect 3960 6610 4310 6620
rect 4320 6610 4350 6620
rect 4370 6610 4380 6620
rect 2220 6600 2370 6610
rect 2440 6600 2510 6610
rect 3680 6600 3710 6610
rect 3800 6600 3890 6610
rect 3940 6600 4360 6610
rect 2210 6590 2340 6600
rect 3670 6590 3690 6600
rect 3790 6590 3870 6600
rect 2220 6580 2330 6590
rect 3770 6580 3850 6590
rect 3900 6580 3920 6590
rect 3930 6580 4370 6600
rect 4410 6590 4420 6600
rect 2230 6570 2310 6580
rect 3900 6570 4380 6580
rect 2240 6560 2300 6570
rect 3890 6560 4360 6570
rect 2240 6540 2290 6560
rect 3880 6550 4340 6560
rect 3790 6540 3820 6550
rect 3840 6540 3890 6550
rect 3950 6540 4350 6550
rect 2230 6530 2270 6540
rect 3760 6530 3900 6540
rect 3970 6530 4360 6540
rect 2240 6520 2260 6530
rect 3759 6520 3960 6530
rect 4000 6520 4360 6530
rect 3720 6519 3738 6520
rect 3720 6510 3750 6519
rect 3760 6510 3980 6520
rect 4010 6510 4370 6520
rect 2240 6500 2250 6510
rect 3730 6500 3740 6510
rect 3790 6500 4390 6510
rect 3810 6490 4390 6500
rect 3800 6470 3810 6480
rect 3830 6470 4340 6490
rect 4362 6480 4410 6490
rect 3750 6460 3920 6470
rect 3940 6460 4340 6470
rect 4350 6465 4386 6480
rect 4430 6470 4450 6490
rect 4350 6460 4380 6465
rect 3760 6450 4010 6460
rect 4020 6450 4380 6460
rect 4480 6450 4500 6480
rect 3730 6440 3740 6450
rect 3770 6440 4310 6450
rect 4320 6440 4380 6450
rect 4510 6440 4530 6450
rect 3770 6430 4300 6440
rect 4320 6430 4390 6440
rect 4510 6430 4540 6440
rect 3780 6420 4390 6430
rect 3790 6410 4320 6420
rect 3700 6400 3710 6410
rect 3730 6400 3840 6410
rect 3760 6390 3840 6400
rect 3870 6390 4270 6410
rect 4290 6400 4330 6410
rect 4340 6400 4390 6420
rect 4320 6390 4400 6400
rect 3770 6380 3860 6390
rect 3870 6380 4280 6390
rect 4330 6380 4350 6390
rect 4390 6380 4420 6390
rect 3790 6360 4290 6380
rect 4440 6369 4461 6381
rect 4450 6360 4460 6369
rect 3800 6350 4300 6360
rect 4370 6350 4390 6360
rect 4450 6350 4470 6360
rect 2180 6340 2190 6350
rect 3800 6340 4280 6350
rect 4370 6340 4400 6350
rect 3800 6330 3830 6340
rect 3840 6330 4260 6340
rect 4270 6330 4290 6340
rect 3800 6320 3820 6330
rect 3860 6320 4250 6330
rect 4280 6320 4290 6330
rect 4380 6320 4400 6340
rect 4450 6330 4490 6350
rect 4470 6320 4490 6330
rect 3810 6310 3830 6320
rect 3870 6310 4250 6320
rect 3820 6300 3840 6310
rect 3870 6300 4260 6310
rect 4310 6300 4320 6310
rect 4440 6300 4450 6310
rect 3740 6290 3750 6300
rect 3830 6290 3850 6300
rect 3880 6290 4040 6300
rect 3830 6270 3860 6290
rect 3890 6280 4040 6290
rect 4050 6280 4060 6290
rect 4070 6280 4270 6300
rect 3910 6270 4060 6280
rect 4080 6270 4270 6280
rect 3510 6250 3520 6270
rect 3770 6260 3780 6270
rect 3810 6260 3870 6270
rect 3920 6260 4070 6270
rect 4090 6260 4270 6270
rect 4420 6260 4430 6280
rect 3770 6250 3790 6260
rect 3780 6240 3790 6250
rect 3820 6250 3880 6260
rect 3910 6250 3950 6260
rect 3980 6250 4040 6260
rect 4050 6250 4280 6260
rect 3820 6240 3890 6250
rect 3900 6240 3950 6250
rect 3620 6210 3630 6220
rect 3750 6219 3760 6240
rect 3820 6230 3880 6240
rect 3900 6230 3910 6240
rect 3810 6220 3880 6230
rect 3940 6220 3960 6240
rect 3990 6230 4000 6250
rect 4010 6240 4040 6250
rect 4060 6240 4090 6250
rect 4020 6231 4040 6240
rect 4020 6220 4050 6231
rect 4070 6230 4090 6240
rect 4110 6240 4290 6250
rect 4110 6230 4300 6240
rect 4070 6220 4100 6230
rect 4120 6220 4200 6230
rect 4220 6220 4300 6230
rect 4350 6220 4360 6250
rect 4430 6240 4440 6250
rect 3750 6210 3771 6219
rect 3790 6210 3890 6220
rect 3620 6200 3640 6210
rect 3760 6200 3890 6210
rect 3930 6200 3960 6220
rect 4029 6219 4050 6220
rect 4040 6210 4050 6219
rect 4080 6210 4150 6220
rect 4030 6200 4150 6210
rect 4170 6210 4210 6220
rect 4221 6210 4310 6220
rect 4170 6200 4230 6210
rect 4240 6200 4310 6210
rect 3750 6190 3780 6200
rect 3800 6190 3900 6200
rect 3930 6190 3970 6200
rect 4030 6190 4320 6200
rect 4450 6190 4460 6198
rect 3640 6189 3650 6190
rect 3639 6177 3660 6189
rect 3760 6180 3780 6190
rect 3790 6180 3820 6190
rect 3650 6170 3660 6177
rect 3590 6150 3600 6160
rect 3650 6150 3670 6170
rect 3700 6150 3730 6170
rect 3480 6140 3490 6150
rect 3590 6140 3610 6150
rect 3590 6130 3620 6140
rect 3660 6130 3680 6150
rect 3520 6120 3530 6130
rect 3580 6120 3630 6130
rect 3650 6120 3680 6130
rect 3710 6130 3730 6150
rect 3750 6160 3820 6180
rect 3840 6170 3900 6190
rect 3940 6180 3980 6190
rect 4030 6180 4120 6190
rect 4130 6180 4180 6190
rect 4200 6180 4320 6190
rect 3940 6170 3990 6180
rect 4020 6170 4120 6180
rect 4140 6170 4180 6180
rect 3840 6160 3910 6170
rect 3940 6160 4000 6170
rect 4020 6160 4060 6170
rect 3750 6140 3830 6160
rect 3840 6150 3920 6160
rect 3940 6150 4010 6160
rect 4035 6159 4056 6160
rect 4040 6150 4050 6159
rect 4070 6150 4110 6170
rect 3740 6130 3830 6140
rect 3850 6140 3930 6150
rect 3940 6140 4020 6150
rect 4040 6140 4110 6150
rect 3850 6130 4030 6140
rect 4050 6130 4110 6140
rect 4150 6160 4180 6170
rect 4210 6170 4320 6180
rect 4440 6170 4480 6190
rect 4210 6160 4310 6170
rect 4150 6140 4190 6160
rect 4230 6150 4310 6160
rect 4360 6160 4370 6170
rect 4430 6160 4480 6170
rect 4230 6140 4320 6150
rect 4330 6140 4340 6150
rect 4360 6140 4380 6160
rect 4430 6150 4470 6160
rect 4430 6140 4460 6150
rect 4150 6130 4160 6140
rect 4180 6130 4200 6140
rect 4240 6130 4340 6140
rect 3710 6120 3830 6130
rect 3860 6120 4040 6130
rect 4060 6120 4120 6130
rect 4190 6120 4220 6130
rect 4250 6120 4350 6130
rect 3430 6110 3450 6120
rect 3510 6110 3540 6120
rect 3560 6110 3570 6120
rect 3580 6110 3840 6120
rect 3860 6110 4000 6120
rect 4010 6110 4040 6120
rect 4070 6110 4140 6120
rect 4200 6110 4220 6120
rect 4260 6110 4350 6120
rect 4370 6120 4380 6140
rect 4440 6130 4470 6140
rect 3490 6100 3500 6110
rect 3520 6100 3680 6110
rect 3700 6100 4150 6110
rect 4180 6100 4230 6110
rect 4260 6102 4360 6110
rect 3520 6090 3690 6100
rect 3710 6090 4160 6100
rect 4180 6090 4240 6100
rect 4272 6090 4360 6102
rect 3510 6080 3570 6090
rect 3510 6070 3520 6080
rect 3500 6060 3520 6070
rect 3540 6070 3570 6080
rect 3580 6070 3690 6090
rect 3720 6080 3890 6090
rect 3730 6070 3890 6080
rect 3900 6070 4160 6090
rect 3540 6060 3700 6070
rect 3730 6060 4160 6070
rect 4190 6078 4260 6090
rect 4281 6080 4360 6090
rect 4370 6090 4390 6120
rect 4450 6110 4470 6130
rect 4450 6100 4480 6110
rect 4370 6080 4400 6090
rect 4190 6060 4270 6078
rect 4300 6060 4400 6080
rect 3500 6050 3710 6060
rect 3720 6050 4020 6060
rect 4050 6050 4170 6060
rect 4190 6050 4420 6060
rect 2730 6040 3030 6050
rect 3500 6040 4030 6050
rect 4040 6040 4430 6050
rect 2670 6030 3090 6040
rect 3490 6030 3650 6040
rect 3660 6030 3870 6040
rect 2570 6020 3140 6030
rect 3550 6020 3640 6030
rect 3690 6020 3860 6030
rect 2530 6010 3170 6020
rect 3560 6010 3640 6020
rect 3660 6010 3860 6020
rect 3890 6020 4430 6040
rect 3890 6010 4450 6020
rect 2260 6000 2280 6010
rect 2500 6000 3210 6010
rect 3570 6000 3650 6010
rect 3660 6000 3840 6010
rect 3900 6000 4450 6010
rect 2240 5990 2330 6000
rect 2490 5990 3050 6000
rect 3120 5990 3250 6000
rect 3570 5990 3670 6000
rect 2190 5980 2330 5990
rect 2470 5980 3050 5990
rect 3140 5980 3290 5990
rect 3550 5980 3670 5990
rect 3700 5990 3840 6000
rect 3910 5990 4430 6000
rect 3700 5980 3870 5990
rect 3900 5980 4420 5990
rect 2130 5970 2350 5980
rect 2470 5970 3060 5980
rect 3130 5970 3360 5980
rect 3560 5970 4100 5980
rect 4120 5970 4180 5980
rect 4200 5970 4420 5980
rect 2040 5960 2350 5970
rect 1980 5950 2350 5960
rect 2480 5960 3080 5970
rect 3090 5960 3410 5970
rect 3570 5960 4420 5970
rect 2480 5950 3450 5960
rect 3570 5950 3790 5960
rect 3807 5952 3980 5960
rect 3807 5950 3960 5952
rect 3990 5950 4130 5960
rect 4140 5950 4420 5960
rect 1940 5940 2340 5950
rect 1920 5930 2340 5940
rect 2480 5940 3530 5950
rect 3560 5940 3831 5950
rect 2480 5930 3730 5940
rect 3770 5930 3840 5940
rect 3860 5930 3960 5950
rect 4020 5940 4410 5950
rect 3970 5930 3990 5940
rect 4030 5930 4410 5940
rect 1900 5920 2340 5930
rect 2390 5920 2400 5930
rect 2440 5920 2450 5930
rect 2470 5920 3170 5930
rect 3270 5920 3740 5930
rect 3770 5920 3780 5930
rect 3790 5920 3910 5930
rect 3930 5920 4010 5930
rect 4050 5920 4250 5930
rect 4260 5920 4410 5930
rect 1880 5910 2350 5920
rect 2390 5910 3150 5920
rect 3340 5910 3750 5920
rect 3760 5910 3780 5920
rect 3800 5910 3920 5920
rect 3940 5910 4010 5920
rect 4060 5910 4430 5920
rect 1850 5900 3130 5910
rect 3430 5900 3840 5910
rect 3870 5900 4020 5910
rect 1830 5890 2420 5900
rect 2430 5890 3120 5900
rect 3500 5890 4030 5900
rect 4070 5890 4410 5910
rect 4420 5900 4430 5910
rect 1820 5880 2380 5890
rect 2440 5880 3110 5890
rect 3560 5880 4040 5890
rect 1800 5870 2370 5880
rect 1790 5860 2370 5870
rect 1770 5850 2370 5860
rect 1770 5840 1790 5850
rect 1820 5840 2370 5850
rect 1770 5830 1780 5840
rect 1820 5820 2300 5840
rect 1810 5810 2300 5820
rect 2310 5810 2370 5840
rect 2460 5870 2520 5880
rect 2530 5870 3110 5880
rect 3610 5870 4040 5880
rect 4080 5880 4410 5890
rect 4420 5880 4430 5890
rect 4080 5870 4430 5880
rect 2460 5860 3100 5870
rect 3660 5860 4420 5870
rect 2460 5850 3070 5860
rect 3680 5859 4410 5860
rect 3680 5850 3940 5859
rect 3960 5850 4410 5859
rect 2460 5810 2520 5850
rect 2530 5810 3060 5850
rect 3690 5840 3950 5850
rect 3970 5840 4410 5850
rect 3690 5830 3800 5840
rect 3810 5830 3960 5840
rect 3980 5830 4030 5840
rect 4040 5830 4400 5840
rect 3690 5820 3970 5830
rect 3990 5820 4400 5830
rect 3650 5810 3660 5820
rect 3690 5810 3980 5820
rect 4000 5810 4400 5820
rect 1790 5800 2360 5810
rect 1770 5780 2360 5800
rect 2470 5780 2520 5810
rect 1770 5770 2350 5780
rect 1800 5760 2350 5770
rect 2480 5760 2520 5780
rect 2540 5800 3060 5810
rect 3590 5800 3990 5810
rect 4000 5800 4050 5810
rect 4140 5800 4400 5810
rect 1810 5750 2340 5760
rect 1820 5740 2340 5750
rect 2480 5740 2530 5760
rect 1820 5730 1900 5740
rect 1910 5730 2310 5740
rect 2320 5730 2330 5740
rect 1820 5720 2310 5730
rect 1850 5710 2310 5720
rect 2490 5720 2530 5740
rect 2540 5730 3070 5800
rect 3540 5790 4020 5800
rect 4160 5790 4390 5800
rect 3530 5770 4000 5790
rect 4180 5780 4390 5790
rect 4190 5770 4390 5780
rect 3530 5760 3990 5770
rect 4200 5760 4380 5770
rect 3540 5750 3630 5760
rect 3670 5750 3970 5760
rect 4210 5750 4380 5760
rect 3560 5740 3570 5750
rect 3690 5740 3830 5750
rect 3850 5740 3930 5750
rect 4220 5740 4380 5750
rect 3700 5730 3810 5740
rect 3850 5730 3880 5740
rect 3900 5730 3930 5740
rect 2490 5710 2540 5720
rect 1870 5680 2300 5710
rect 2500 5700 2540 5710
rect 2550 5700 3070 5730
rect 2500 5690 2530 5700
rect 2560 5690 3070 5700
rect 3730 5710 3800 5730
rect 3860 5720 3870 5730
rect 4230 5720 4380 5740
rect 4120 5710 4130 5720
rect 4240 5710 4380 5720
rect 1880 5670 1890 5680
rect 1900 5670 2300 5680
rect 2560 5670 3060 5690
rect 3730 5680 3760 5710
rect 3770 5700 3800 5710
rect 4150 5700 4160 5710
rect 4250 5700 4380 5710
rect 3770 5690 3790 5700
rect 4010 5690 4040 5700
rect 4150 5690 4180 5700
rect 4260 5690 4380 5700
rect 3710 5670 3760 5680
rect 4000 5670 4030 5690
rect 4160 5680 4190 5690
rect 4260 5680 4370 5690
rect 4170 5670 4200 5680
rect 4270 5670 4370 5680
rect 1880 5650 2310 5670
rect 1880 5610 2300 5650
rect 2540 5640 2550 5649
rect 2540 5630 2560 5640
rect 2570 5630 3060 5670
rect 3100 5660 3120 5670
rect 3710 5660 3730 5670
rect 3620 5650 3640 5660
rect 3600 5640 3640 5650
rect 3700 5650 3730 5660
rect 3700 5640 3710 5650
rect 3990 5640 4030 5670
rect 4180 5660 4210 5670
rect 4160 5650 4220 5660
rect 4270 5650 4360 5670
rect 4200 5640 4220 5650
rect 3600 5630 3630 5640
rect 3690 5630 3710 5640
rect 4180 5630 4220 5640
rect 4280 5640 4310 5650
rect 4320 5640 4360 5650
rect 2550 5620 2560 5630
rect 2580 5610 3060 5630
rect 3610 5620 3630 5630
rect 3660 5620 3680 5630
rect 3650 5610 3680 5620
rect 4190 5620 4230 5630
rect 4280 5620 4300 5640
rect 4340 5630 4350 5640
rect 1880 5590 2290 5610
rect 2590 5590 3050 5610
rect 3650 5600 3670 5610
rect 1880 5560 2280 5590
rect 2600 5580 3040 5590
rect 2610 5570 3040 5580
rect 3960 5580 3980 5590
rect 4190 5580 4220 5620
rect 3960 5570 4000 5580
rect 2610 5560 3030 5570
rect 1890 5530 2270 5560
rect 2620 5550 3030 5560
rect 3950 5560 4020 5570
rect 4200 5560 4220 5580
rect 4280 5610 4310 5620
rect 4280 5600 4340 5610
rect 4280 5590 4310 5600
rect 4320 5590 4330 5600
rect 4280 5560 4330 5590
rect 3950 5550 4030 5560
rect 4200 5550 4230 5560
rect 2630 5530 3020 5550
rect 3950 5540 4050 5550
rect 3960 5530 4050 5540
rect 4200 5530 4220 5550
rect 4280 5540 4320 5560
rect 1900 5520 2270 5530
rect 2650 5520 3010 5530
rect 3960 5520 4060 5530
rect 1900 5500 2260 5520
rect 2660 5510 3000 5520
rect 2670 5500 2990 5510
rect 1910 5480 2250 5500
rect 2570 5490 2600 5500
rect 2690 5490 2970 5500
rect 3960 5490 4000 5520
rect 4020 5510 4040 5520
rect 4200 5510 4210 5530
rect 4280 5510 4290 5540
rect 4300 5530 4320 5540
rect 4020 5490 4030 5510
rect 4270 5500 4290 5510
rect 2520 5480 2530 5490
rect 2560 5480 2610 5490
rect 2710 5480 2950 5490
rect 3970 5480 3990 5490
rect 4270 5480 4300 5500
rect 1920 5470 2250 5480
rect 2560 5470 2620 5480
rect 2710 5470 2930 5480
rect 4260 5470 4280 5480
rect 1930 5450 2240 5470
rect 2560 5460 2640 5470
rect 2690 5460 2880 5470
rect 4260 5460 4270 5470
rect 4290 5460 4300 5480
rect 2570 5450 2650 5460
rect 2680 5450 2740 5460
rect 4250 5450 4270 5460
rect 1940 5440 2230 5450
rect 1950 5430 2220 5440
rect 2580 5430 2730 5450
rect 3910 5430 3920 5440
rect 1960 5420 2210 5430
rect 2580 5420 2690 5430
rect 2700 5420 2730 5430
rect 3930 5420 3950 5430
rect 4240 5420 4270 5450
rect 1970 5410 2210 5420
rect 2590 5410 2690 5420
rect 3940 5410 3950 5420
rect 4080 5410 4100 5420
rect 4230 5410 4260 5420
rect 1990 5400 2200 5410
rect 2600 5400 2710 5410
rect 2030 5390 2110 5400
rect 2170 5390 2200 5400
rect 2610 5390 2710 5400
rect 4220 5390 4260 5410
rect 2180 5380 2190 5390
rect 2600 5380 2720 5390
rect 2610 5370 2730 5380
rect 4210 5370 4250 5390
rect 2610 5360 2740 5370
rect 2240 5350 2260 5360
rect 2610 5350 2750 5360
rect 4200 5350 4250 5370
rect 2240 5340 2270 5350
rect 2600 5340 2760 5350
rect 4190 5340 4240 5350
rect 2250 5330 2290 5340
rect 2600 5330 2770 5340
rect 2250 5320 2300 5330
rect 2420 5320 2530 5330
rect 2590 5320 2770 5330
rect 4180 5320 4240 5340
rect 2260 5310 2310 5320
rect 2380 5310 2550 5320
rect 2580 5310 2790 5320
rect 4170 5310 4230 5320
rect 2260 5300 2330 5310
rect 2350 5300 2790 5310
rect 4160 5300 4230 5310
rect 2260 5290 2340 5300
rect 2350 5290 2800 5300
rect 4150 5290 4230 5300
rect 2260 5280 2800 5290
rect 4140 5280 4220 5290
rect 2230 5270 2610 5280
rect 2640 5270 2800 5280
rect 4130 5270 4220 5280
rect 2230 5260 2590 5270
rect 2640 5260 2810 5270
rect 4120 5260 4210 5270
rect 2220 5250 2370 5260
rect 2380 5250 2590 5260
rect 2660 5250 2810 5260
rect 3850 5250 3890 5260
rect 4110 5250 4210 5260
rect 2220 5240 2610 5250
rect 2690 5241 2810 5250
rect 2712 5240 2810 5241
rect 4100 5240 4200 5250
rect 2220 5220 2320 5240
rect 2330 5230 2610 5240
rect 2720 5230 2810 5240
rect 4090 5230 4200 5240
rect 2090 5200 2110 5220
rect 2220 5210 2310 5220
rect 2350 5210 2530 5230
rect 2550 5220 2610 5230
rect 2712 5229 2810 5230
rect 2700 5220 2810 5229
rect 2840 5220 2850 5230
rect 4090 5220 4190 5230
rect 2540 5210 2600 5220
rect 2730 5210 2820 5220
rect 2220 5200 2290 5210
rect 2210 5190 2290 5200
rect 2350 5200 2590 5210
rect 2740 5200 2830 5210
rect 3780 5200 3810 5210
rect 2350 5190 2580 5200
rect 2750 5190 2840 5200
rect 3770 5190 3810 5200
rect 4080 5190 4180 5220
rect 2210 5180 2280 5190
rect 2080 5160 2130 5180
rect 2090 5150 2130 5160
rect 2200 5170 2270 5180
rect 2370 5170 2580 5190
rect 2760 5180 2850 5190
rect 2640 5170 2660 5180
rect 2790 5170 2840 5180
rect 3770 5170 3800 5190
rect 4070 5170 4170 5190
rect 2200 5160 2260 5170
rect 2350 5160 2480 5170
rect 2520 5160 2530 5170
rect 2540 5160 2580 5170
rect 3770 5160 3790 5170
rect 4070 5160 4160 5170
rect 2200 5150 2250 5160
rect 2080 5140 2130 5150
rect 2210 5140 2250 5150
rect 2350 5150 2470 5160
rect 2550 5150 2580 5160
rect 4060 5150 4160 5160
rect 2350 5140 2480 5150
rect 2570 5140 2590 5150
rect 4060 5140 4150 5150
rect 2080 5130 2140 5140
rect 2070 5120 2140 5130
rect 2200 5130 2240 5140
rect 2200 5120 2230 5130
rect 2350 5120 2460 5140
rect 2040 5100 2050 5120
rect 2060 5100 2150 5120
rect 2200 5110 2220 5120
rect 2340 5110 2460 5120
rect 4050 5120 4140 5140
rect 4050 5110 4110 5120
rect 4120 5110 4130 5120
rect 2070 5070 2150 5100
rect 2340 5100 2450 5110
rect 2340 5090 2430 5100
rect 4040 5090 4110 5110
rect 2380 5080 2410 5090
rect 2080 5060 2150 5070
rect 4030 5070 4110 5090
rect 4030 5060 4100 5070
rect 2080 5030 2160 5060
rect 2450 5050 2520 5060
rect 4030 5050 4090 5060
rect 2320 5040 2350 5050
rect 2430 5040 2560 5050
rect 2320 5030 2390 5040
rect 2410 5030 2600 5040
rect 4020 5030 4090 5050
rect 2090 5010 2160 5030
rect 2310 5020 2630 5030
rect 2300 5010 2660 5020
rect 4020 5010 4070 5030
rect 2100 5000 2160 5010
rect 2301 5000 2690 5010
rect 2120 4990 2150 5000
rect 2301 4990 2700 5000
rect 2720 4990 2790 5000
rect 4010 4990 4060 5010
rect 2301 4989 2830 4990
rect 2280 4980 2290 4986
rect 2300 4980 2830 4989
rect 2280 4970 2850 4980
rect 4010 4970 4050 4990
rect 2220 4960 2230 4970
rect 2270 4960 2860 4970
rect 2210 4950 2240 4960
rect 2270 4950 2870 4960
rect 4000 4950 4040 4970
rect 2210 4940 2530 4950
rect 2600 4940 2620 4950
rect 2630 4940 2890 4950
rect 2210 4930 2480 4940
rect 2670 4930 2690 4940
rect 2720 4930 2890 4940
rect 2210 4920 2440 4930
rect 2750 4920 2900 4930
rect 4000 4920 4030 4950
rect 2210 4910 2322 4920
rect 2352 4910 2430 4920
rect 2810 4910 2910 4920
rect 2210 4900 2320 4910
rect 2370 4900 2400 4910
rect 2830 4900 2890 4910
rect 2900 4900 2910 4910
rect 2210 4880 2310 4900
rect 2370 4890 2380 4900
rect 2360 4880 2380 4890
rect 2850 4890 2880 4900
rect 2900 4890 2920 4900
rect 3990 4890 4020 4920
rect 2850 4880 2930 4890
rect 3990 4880 4010 4890
rect 2210 4870 2300 4880
rect 2220 4860 2280 4870
rect 2360 4860 2370 4880
rect 2500 4870 2510 4880
rect 2870 4870 2930 4880
rect 2390 4860 2430 4870
rect 2880 4860 2930 4870
rect 2220 4850 2260 4860
rect 2360 4850 2450 4860
rect 2890 4850 2930 4860
rect 2230 4820 2260 4850
rect 2330 4840 2460 4850
rect 2910 4840 2930 4850
rect 3980 4870 4010 4880
rect 3980 4850 4000 4870
rect 2320 4830 2460 4840
rect 3980 4830 3990 4850
rect 2330 4820 2460 4830
rect 2240 4810 2250 4820
rect 2340 4810 2480 4820
rect 2330 4800 2510 4810
rect 3970 4800 3980 4820
rect 2330 4780 2530 4800
rect 2320 4770 2540 4780
rect 2570 4770 2600 4780
rect 2330 4760 2650 4770
rect 2090 4750 2110 4760
rect 2130 4750 2140 4760
rect 2330 4750 2670 4760
rect 2340 4730 2700 4750
rect 2000 4710 2070 4730
rect 2330 4720 2710 4730
rect 2330 4710 2720 4720
rect 2010 4700 2050 4710
rect 2330 4700 2730 4710
rect 1080 4690 1090 4700
rect 2010 4690 2080 4700
rect 2210 4690 2220 4700
rect 2330 4690 2740 4700
rect 1050 4680 1090 4690
rect 1040 4670 1090 4680
rect 2020 4670 2090 4690
rect 2340 4680 2740 4690
rect 2340 4670 2730 4680
rect 1030 4660 1050 4670
rect 1030 4640 1040 4660
rect 1080 4650 1090 4670
rect 2050 4660 2080 4670
rect 2330 4660 2710 4670
rect 1800 4650 1810 4660
rect 2030 4650 2080 4660
rect 2340 4650 2700 4660
rect 1780 4640 1810 4650
rect 2010 4610 2070 4650
rect 2340 4641 2560 4650
rect 2340 4640 2544 4641
rect 2600 4640 2700 4650
rect 2350 4632 2544 4640
rect 2350 4630 2520 4632
rect 2620 4630 2670 4640
rect 2360 4620 2520 4630
rect 2370 4610 2410 4620
rect 2450 4610 2520 4620
rect 1030 4590 1040 4610
rect 2010 4590 2050 4610
rect 2370 4600 2390 4610
rect 2460 4600 2510 4610
rect 2530 4600 2540 4620
rect 2010 4580 2070 4590
rect 2010 4570 2080 4580
rect 2450 4570 2520 4600
rect 5800 4570 5810 4590
rect 1940 4560 1990 4570
rect 2000 4560 2090 4570
rect 2280 4560 2310 4570
rect 1930 4550 2090 4560
rect 2290 4550 2310 4560
rect 1920 4540 2090 4550
rect 2300 4540 2320 4550
rect 2450 4540 2530 4570
rect 1920 4530 1990 4540
rect 2010 4530 2120 4540
rect 2210 4530 2250 4540
rect 2450 4530 2540 4540
rect 1920 4510 1970 4530
rect 2020 4521 2130 4530
rect 2020 4520 2109 4521
rect 2440 4520 2550 4530
rect 2030 4510 2109 4520
rect 2430 4510 2560 4520
rect 2040 4490 2090 4510
rect 2270 4500 2300 4510
rect 2280 4490 2300 4500
rect 2040 4480 2050 4490
rect 2060 4480 2080 4490
rect 1010 4460 1030 4470
rect 2070 4460 2080 4480
rect 2310 4470 2320 4490
rect 2450 4480 2570 4510
rect 2400 4470 2590 4480
rect 2410 4460 2600 4470
rect 2400 4450 2600 4460
rect 2400 4440 2680 4450
rect 1010 4420 1030 4440
rect 2400 4430 2690 4440
rect 2710 4430 2720 4440
rect 2320 4420 2340 4430
rect 2400 4420 2750 4430
rect 2260 4419 2271 4420
rect 2260 4410 2290 4419
rect 2280 4400 2290 4410
rect 2400 4410 2760 4420
rect 2400 4400 2790 4410
rect 2400 4390 2820 4400
rect 2400 4380 2830 4390
rect 2410 4360 2850 4380
rect 2880 4370 2910 4380
rect 2890 4360 2910 4370
rect 2380 4350 2400 4360
rect 2420 4350 2860 4360
rect 3240 4350 3250 4360
rect 2410 4340 2870 4350
rect 2900 4340 2910 4350
rect 3050 4340 3080 4350
rect 3090 4340 3150 4350
rect 3210 4340 3230 4350
rect 3960 4340 3970 4350
rect 2340 4330 2350 4340
rect 2410 4330 2850 4340
rect 2880 4330 2950 4340
rect 3010 4330 3250 4340
rect 2280 4310 2290 4330
rect 2340 4320 2360 4330
rect 2450 4320 2840 4330
rect 2480 4310 2840 4320
rect 2870 4320 2970 4330
rect 2990 4320 3250 4330
rect 3950 4320 3980 4340
rect 2870 4310 3220 4320
rect 3950 4310 3960 4320
rect 2270 4300 2290 4310
rect 2310 4300 2330 4310
rect 2350 4300 2370 4310
rect 2490 4300 3220 4310
rect 2260 4290 2400 4300
rect 2480 4290 3230 4300
rect 3940 4290 3960 4310
rect 3990 4300 4010 4310
rect 4000 4290 4010 4300
rect 2250 4280 2420 4290
rect 2250 4270 2330 4280
rect 2360 4270 2420 4280
rect 2470 4270 2680 4290
rect 2700 4280 2760 4290
rect 2770 4280 3230 4290
rect 3950 4280 3970 4290
rect 2230 4260 2280 4270
rect 2310 4260 2430 4270
rect 2460 4260 2680 4270
rect 2710 4260 2780 4280
rect 2800 4270 3250 4280
rect 3950 4270 3990 4280
rect 2810 4260 3270 4270
rect 1890 4250 1900 4260
rect 2190 4250 2290 4260
rect 1970 4230 1980 4250
rect 2100 4240 2290 4250
rect 2090 4230 2290 4240
rect 2300 4250 2420 4260
rect 2450 4250 2680 4260
rect 2730 4250 2780 4260
rect 2300 4240 2700 4250
rect 2740 4240 2790 4250
rect 2820 4240 3280 4260
rect 3960 4250 3990 4270
rect 3970 4240 3990 4250
rect 2300 4230 2710 4240
rect 1920 4220 1980 4230
rect 2080 4220 2200 4230
rect 930 4210 940 4220
rect 1910 4210 1980 4220
rect 2070 4210 2200 4220
rect 2210 4220 2660 4230
rect 2210 4210 2230 4220
rect 2260 4210 2650 4220
rect 2670 4210 2710 4230
rect 2740 4230 2800 4240
rect 2810 4230 3290 4240
rect 3980 4230 3990 4240
rect 2740 4220 2830 4230
rect 2860 4220 3290 4230
rect 3950 4220 3960 4230
rect 2750 4210 2830 4220
rect 550 4200 570 4210
rect 530 4190 570 4200
rect 920 4200 950 4210
rect 1870 4200 1881 4210
rect 1920 4200 1990 4210
rect 2070 4200 2220 4210
rect 2260 4200 2660 4210
rect 2670 4200 2720 4210
rect 2770 4200 2830 4210
rect 2870 4200 3290 4220
rect 540 4180 590 4190
rect 920 4180 960 4200
rect 1890 4190 2000 4200
rect 2060 4190 2740 4200
rect 540 4160 580 4180
rect 930 4170 960 4180
rect 1870 4180 2010 4190
rect 2060 4180 2370 4190
rect 2380 4180 2680 4190
rect 2690 4180 2740 4190
rect 2780 4190 2840 4200
rect 2870 4190 3280 4200
rect 2780 4180 2850 4190
rect 2860 4180 3290 4190
rect 1870 4170 2050 4180
rect 2060 4170 2680 4180
rect 940 4160 980 4170
rect 1870 4160 2680 4170
rect 530 4150 590 4160
rect 940 4150 970 4160
rect 1870 4150 2290 4160
rect 2300 4150 2680 4160
rect 520 4100 590 4150
rect 930 4140 960 4150
rect 910 4130 960 4140
rect 1870 4140 2320 4150
rect 2330 4140 2680 4150
rect 2700 4160 2750 4180
rect 2780 4160 2890 4180
rect 2920 4170 3280 4180
rect 3940 4170 3960 4220
rect 3990 4200 4000 4210
rect 2700 4140 2790 4160
rect 2820 4150 2890 4160
rect 1870 4130 2310 4140
rect 2330 4130 2710 4140
rect 2730 4130 2790 4140
rect 920 4122 960 4130
rect 942 4110 960 4122
rect 1900 4120 2300 4130
rect 1910 4110 2100 4120
rect 2110 4110 2280 4120
rect 530 4080 590 4100
rect 1930 4090 2060 4110
rect 2150 4100 2250 4110
rect 2320 4100 2710 4130
rect 2740 4120 2790 4130
rect 2830 4140 2890 4150
rect 2930 4160 3270 4170
rect 2930 4150 3260 4160
rect 3940 4150 3970 4170
rect 2930 4140 3270 4150
rect 3940 4140 3980 4150
rect 2830 4130 3290 4140
rect 2740 4110 2800 4120
rect 2830 4110 2950 4130
rect 2990 4110 3290 4130
rect 2740 4100 2850 4110
rect 2880 4100 2950 4110
rect 3000 4100 3310 4110
rect 3940 4100 3990 4140
rect 2160 4090 2210 4100
rect 2220 4090 2260 4100
rect 2310 4090 2720 4100
rect 2750 4092 2850 4100
rect 2769 4090 2850 4092
rect 1940 4080 2050 4090
rect 2170 4080 2210 4090
rect 2240 4080 2260 4090
rect 2300 4080 2730 4090
rect 2780 4080 2850 4090
rect 2890 4090 2960 4100
rect 2990 4090 3310 4100
rect 2890 4080 2970 4090
rect 2990 4080 3020 4090
rect 3040 4080 3310 4090
rect 3930 4090 3980 4100
rect 3930 4080 3970 4090
rect 520 4070 590 4080
rect 1950 4070 2040 4080
rect 2240 4070 2250 4080
rect 2300 4070 2750 4080
rect 560 4060 590 4070
rect 2020 4060 2040 4070
rect 2170 4060 2180 4070
rect 2290 4060 2750 4070
rect 2790 4070 2850 4080
rect 2900 4070 3020 4080
rect 3060 4070 3310 4080
rect 2790 4060 2860 4070
rect 2890 4060 3010 4070
rect 3060 4060 3150 4070
rect 3160 4060 3310 4070
rect 3920 4060 3960 4080
rect 2170 4040 2200 4060
rect 2210 4040 2220 4060
rect 2290 4050 2760 4060
rect 2270 4040 2760 4050
rect 2800 4041 2910 4060
rect 2940 4050 3020 4060
rect 2820 4040 2910 4041
rect 2950 4040 3020 4050
rect 3070 4050 3320 4060
rect 3910 4050 3950 4060
rect 3070 4040 3330 4050
rect 3910 4040 3940 4050
rect 2170 4030 2180 4040
rect 2270 4030 2780 4040
rect 850 4020 860 4030
rect 920 4020 940 4030
rect 2260 4029 2793 4030
rect 2260 4020 2800 4029
rect 2840 4020 2910 4040
rect 2960 4030 3030 4040
rect 3060 4030 3100 4040
rect 3110 4030 3340 4040
rect 3900 4030 3930 4040
rect 2960 4020 3090 4030
rect 890 4010 900 4020
rect 880 4000 900 4010
rect 920 4010 950 4020
rect 2250 4010 2800 4020
rect 2850 4010 2920 4020
rect 2950 4010 3080 4020
rect 3130 4010 3210 4030
rect 3250 4020 3339 4030
rect 3890 4020 3920 4030
rect 4180 4020 4190 4030
rect 3250 4010 3310 4020
rect 3330 4010 3340 4020
rect 3890 4010 3910 4020
rect 920 4000 960 4010
rect 2240 4000 2810 4010
rect 910 3990 960 4000
rect 2180 3990 2190 4000
rect 2230 3990 2810 4000
rect 2860 4000 2930 4010
rect 2940 4000 2970 4010
rect 3010 4000 3080 4010
rect 3140 4000 3220 4010
rect 3250 4000 3340 4010
rect 3880 4000 3900 4010
rect 2860 3990 2970 4000
rect 910 3980 970 3990
rect 2090 3980 2110 3990
rect 2170 3980 2190 3990
rect 2220 3980 2820 3990
rect 2850 3980 2870 3990
rect 2890 3980 2970 3990
rect 3020 3990 3090 4000
rect 3140 3990 3300 4000
rect 3310 3990 3350 4000
rect 3880 3990 3890 4000
rect 3020 3980 3100 3990
rect 3130 3980 3280 3990
rect 3330 3980 3370 3990
rect 910 3970 990 3980
rect 2210 3970 2860 3980
rect 900 3960 1000 3970
rect 2070 3960 2090 3970
rect 2130 3960 2860 3970
rect 2910 3970 2970 3980
rect 3030 3970 3150 3980
rect 3200 3970 3280 3980
rect 3350 3970 3390 3980
rect 5560 3970 5570 3990
rect 2910 3960 2980 3970
rect 3010 3960 3150 3970
rect 900 3950 1010 3960
rect 2050 3950 2780 3960
rect 2800 3950 2870 3960
rect 910 3930 1010 3950
rect 2010 3940 2780 3950
rect 1980 3930 2780 3940
rect 2810 3940 2870 3950
rect 2920 3950 3040 3960
rect 3070 3950 3150 3960
rect 2920 3940 3030 3950
rect 2810 3930 2890 3940
rect 2920 3939 2930 3940
rect 2960 3930 3030 3940
rect 3090 3940 3150 3950
rect 3210 3950 3280 3970
rect 3360 3960 3390 3970
rect 3210 3940 3279 3950
rect 3090 3930 3160 3940
rect 3255 3939 3280 3940
rect 3270 3930 3280 3939
rect 900 3920 1010 3930
rect 1940 3920 2790 3930
rect 2820 3920 2920 3930
rect 890 3910 1020 3920
rect 1870 3910 2920 3920
rect 2970 3920 3040 3930
rect 3100 3920 3190 3930
rect 3290 3920 3330 3930
rect 2970 3910 3050 3920
rect 3100 3910 3200 3920
rect 890 3900 1010 3910
rect 1820 3900 2830 3910
rect 2860 3900 2930 3910
rect 850 3880 870 3890
rect 880 3880 1010 3900
rect 1790 3890 2830 3900
rect 1760 3880 2830 3890
rect 850 3870 1010 3880
rect 1730 3870 2830 3880
rect 2870 3890 2930 3900
rect 2980 3900 3060 3910
rect 3080 3900 3090 3910
rect 3140 3900 3210 3910
rect 3290 3900 3340 3920
rect 3440 3910 3450 3940
rect 4060 3930 4080 3950
rect 5930 3940 5940 3960
rect 4060 3920 4090 3930
rect 5410 3920 5420 3930
rect 4060 3900 4100 3920
rect 5570 3910 5590 3920
rect 2980 3890 3100 3900
rect 3150 3890 3220 3900
rect 3300 3890 3350 3900
rect 2870 3880 2950 3890
rect 2970 3880 2990 3890
rect 3020 3880 3100 3890
rect 2870 3870 2990 3880
rect 900 3860 1010 3870
rect 1700 3860 2850 3870
rect 2860 3860 2990 3870
rect 850 3830 870 3860
rect 900 3850 1020 3860
rect 1680 3850 2890 3860
rect 2920 3850 2990 3860
rect 910 3840 1030 3850
rect 1650 3840 2880 3850
rect 2930 3840 2990 3850
rect 3040 3870 3100 3880
rect 3170 3880 3220 3890
rect 3320 3880 3330 3890
rect 4070 3880 4100 3900
rect 5560 3900 5600 3910
rect 5560 3890 5590 3900
rect 5850 3890 5880 3900
rect 5840 3880 5880 3890
rect 3170 3870 3230 3880
rect 3370 3870 3400 3880
rect 4060 3870 4100 3880
rect 5829 3870 5880 3880
rect 3040 3850 3110 3870
rect 3190 3860 3240 3870
rect 3360 3860 3410 3870
rect 3220 3850 3280 3860
rect 3040 3840 3150 3850
rect 3230 3840 3290 3850
rect 3370 3840 3410 3860
rect 3510 3860 3520 3870
rect 4060 3860 4110 3870
rect 5480 3860 5490 3870
rect 3510 3850 3530 3860
rect 4060 3840 4130 3860
rect 5480 3850 5500 3860
rect 5480 3840 5530 3850
rect 910 3830 1020 3840
rect 1600 3830 2890 3840
rect 2930 3830 3010 3840
rect 3090 3830 3160 3840
rect 910 3820 1010 3830
rect 1570 3820 2890 3830
rect 2940 3820 3040 3830
rect 3100 3820 3160 3830
rect 3240 3820 3290 3840
rect 4060 3830 4140 3840
rect 4900 3830 4910 3840
rect 4060 3820 4150 3830
rect 4707 3822 4730 3830
rect 4690 3820 4730 3822
rect 4880 3820 4920 3830
rect 5470 3820 5530 3840
rect 910 3810 1000 3820
rect 1550 3810 2900 3820
rect 2930 3810 3050 3820
rect 910 3800 930 3810
rect 1520 3800 2950 3810
rect 920 3790 930 3800
rect 1490 3790 2950 3800
rect 2990 3800 3050 3810
rect 3110 3810 3170 3820
rect 3250 3810 3290 3820
rect 3110 3800 3180 3810
rect 3300 3800 3340 3810
rect 2990 3790 3060 3800
rect 3120 3790 3210 3800
rect 890 3780 910 3790
rect 1460 3780 2940 3790
rect 3000 3780 3070 3790
rect 3150 3780 3220 3790
rect 3300 3780 3360 3800
rect 3440 3790 3480 3820
rect 3580 3810 3590 3820
rect 3720 3810 3740 3820
rect 3580 3800 3600 3810
rect 3720 3800 3770 3810
rect 3710 3790 3780 3800
rect 3450 3780 3470 3790
rect 3600 3780 3620 3790
rect 3680 3780 3790 3790
rect 4060 3780 4160 3820
rect 4680 3810 4740 3820
rect 4670 3800 4740 3810
rect 4880 3810 4940 3820
rect 5470 3810 5490 3820
rect 4670 3780 4750 3800
rect 4880 3780 4930 3810
rect 5330 3800 5340 3810
rect 5450 3800 5510 3810
rect 5330 3790 5360 3800
rect 5440 3790 5510 3800
rect 5670 3790 5690 3800
rect 130 3770 140 3780
rect 880 3770 900 3780
rect 1440 3770 2860 3780
rect 2880 3770 2950 3780
rect 3000 3770 3100 3780
rect 3170 3770 3230 3780
rect 3310 3770 3350 3780
rect 3600 3770 3630 3780
rect 3660 3770 3800 3780
rect 4060 3770 4170 3780
rect 4210 3770 4240 3780
rect 4670 3770 4760 3780
rect 690 3760 710 3770
rect 879 3768 890 3770
rect 670 3750 730 3760
rect 650 3740 740 3750
rect 800 3740 830 3760
rect 860 3740 890 3768
rect 1410 3760 2860 3770
rect 1400 3750 2860 3760
rect 2890 3760 2960 3770
rect 2990 3760 3110 3770
rect 2890 3750 3010 3760
rect 3050 3750 3120 3760
rect 3180 3750 3240 3770
rect 3330 3760 3350 3770
rect 3590 3760 3630 3770
rect 3650 3760 3810 3770
rect 4060 3760 4260 3770
rect 4660 3760 4770 3770
rect 4890 3760 4930 3780
rect 5320 3780 5360 3790
rect 5380 3780 5410 3790
rect 5450 3780 5480 3790
rect 5490 3780 5510 3790
rect 5320 3770 5430 3780
rect 5440 3770 5500 3780
rect 5320 3760 5500 3770
rect 5660 3770 5780 3790
rect 5960 3780 5970 3790
rect 5990 3780 6000 3790
rect 5950 3770 5970 3780
rect 5980 3770 6010 3780
rect 5660 3760 5790 3770
rect 3380 3750 3400 3760
rect 3520 3750 3550 3760
rect 3590 3750 3620 3760
rect 3650 3750 3820 3760
rect 4060 3750 4290 3760
rect 4670 3750 4770 3760
rect 1370 3740 2870 3750
rect 2890 3740 3000 3750
rect 640 3730 780 3740
rect 790 3730 840 3740
rect 860 3730 880 3740
rect 1310 3730 2910 3740
rect 2930 3730 3010 3740
rect 3060 3730 3130 3750
rect 3190 3740 3240 3750
rect 3250 3740 3260 3750
rect 3380 3740 3420 3750
rect 3510 3740 3550 3750
rect 3660 3740 3830 3750
rect 3230 3730 3290 3740
rect 650 3720 870 3730
rect 1290 3720 2910 3730
rect 2940 3720 3010 3730
rect 3070 3720 3150 3730
rect 3240 3720 3300 3730
rect 3380 3720 3430 3740
rect 3520 3730 3550 3740
rect 3680 3730 3830 3740
rect 4060 3740 4300 3750
rect 4670 3740 4760 3750
rect 4870 3740 4940 3760
rect 5310 3750 5500 3760
rect 5640 3750 5650 3760
rect 5660 3750 5810 3760
rect 5940 3750 6010 3770
rect 4060 3730 4340 3740
rect 4660 3730 4750 3740
rect 4890 3730 4930 3740
rect 5300 3730 5510 3750
rect 5640 3740 5810 3750
rect 5970 3740 5990 3750
rect 5640 3730 5800 3740
rect 5970 3730 5980 3740
rect 3680 3720 3840 3730
rect 4060 3720 4350 3730
rect 4670 3720 4750 3730
rect 650 3710 860 3720
rect 1260 3710 2910 3720
rect 660 3700 890 3710
rect 1250 3700 2910 3710
rect 2950 3710 3020 3720
rect 3080 3710 3180 3720
rect 2950 3700 3040 3710
rect 3120 3700 3190 3710
rect 3250 3700 3310 3720
rect 3390 3710 3420 3720
rect 3570 3710 3580 3720
rect 3690 3710 3850 3720
rect 3550 3700 3590 3710
rect 3700 3700 3850 3710
rect 4060 3710 4400 3720
rect 4680 3710 4750 3720
rect 4900 3720 4920 3730
rect 5310 3720 5520 3730
rect 5650 3720 5780 3730
rect 5960 3720 5980 3730
rect 4900 3710 4910 3720
rect 5340 3710 5530 3720
rect 5650 3710 5760 3720
rect 5950 3710 5980 3720
rect 50 3690 60 3700
rect 50 3680 70 3690
rect 660 3680 900 3700
rect 1220 3690 2920 3700
rect 2950 3690 3070 3700
rect 1170 3680 2930 3690
rect 2950 3680 2970 3690
rect 3000 3680 3070 3690
rect 3130 3690 3190 3700
rect 3260 3690 3310 3700
rect 3480 3690 3490 3700
rect 3130 3680 3200 3690
rect 3290 3680 3320 3690
rect 3330 3680 3350 3690
rect 3470 3680 3500 3690
rect 50 3670 60 3680
rect 670 3670 800 3680
rect 820 3670 880 3680
rect 1120 3670 2960 3680
rect 3010 3670 3080 3680
rect 3140 3670 3210 3680
rect 3310 3670 3360 3680
rect 3460 3670 3500 3680
rect 3550 3680 3580 3700
rect 3700 3690 3860 3700
rect 3650 3680 3730 3690
rect 3550 3670 3590 3680
rect 3600 3670 3720 3680
rect 3750 3670 3870 3690
rect 4060 3680 4240 3710
rect 4260 3700 4410 3710
rect 4670 3700 4740 3710
rect 5310 3700 5520 3710
rect 5640 3700 5770 3710
rect 4270 3690 4450 3700
rect 4670 3690 4730 3700
rect 4870 3690 4930 3700
rect 5310 3690 5530 3700
rect 5640 3690 5760 3700
rect 5840 3690 5850 3700
rect 4270 3680 4460 3690
rect 4060 3670 4250 3680
rect 4290 3670 4460 3680
rect 4670 3670 4720 3690
rect 5310 3670 5370 3690
rect 5390 3680 5540 3690
rect 5410 3670 5550 3680
rect 670 3660 680 3670
rect 690 3660 750 3670
rect 770 3660 800 3670
rect 830 3660 880 3670
rect 1110 3660 2960 3670
rect 3020 3660 3080 3670
rect 3150 3660 3240 3670
rect 3320 3660 3370 3670
rect 3460 3660 3490 3670
rect 3560 3660 3680 3670
rect 3690 3660 3720 3670
rect 3770 3660 3801 3670
rect 690 3650 760 3660
rect 790 3650 820 3660
rect 830 3650 940 3660
rect 1090 3650 2970 3660
rect 3020 3650 3090 3660
rect 3180 3650 3250 3660
rect 3320 3650 3380 3660
rect 3550 3651 3720 3660
rect 3550 3650 3732 3651
rect 690 3640 770 3650
rect 700 3630 770 3640
rect 790 3640 920 3650
rect 930 3640 940 3650
rect 1010 3640 2980 3650
rect 3030 3640 3130 3650
rect 3190 3640 3260 3650
rect 3330 3640 3370 3650
rect 3510 3640 3650 3650
rect 3660 3640 3680 3650
rect 3710 3642 3732 3650
rect 3780 3648 3801 3660
rect 3810 3660 3880 3670
rect 4060 3660 4260 3670
rect 3810 3650 3820 3660
rect 3710 3640 3741 3642
rect 3790 3640 3800 3648
rect 3830 3640 3890 3660
rect 4060 3650 4270 3660
rect 4060 3640 4290 3650
rect 4300 3640 4490 3670
rect 4670 3660 4730 3670
rect 5280 3660 5290 3670
rect 4530 3640 4550 3660
rect 790 3630 910 3640
rect 990 3630 2990 3640
rect 3060 3630 3140 3640
rect 3200 3630 3270 3640
rect 3350 3630 3370 3640
rect 3500 3630 3670 3640
rect 3717 3630 3760 3640
rect 3820 3630 3840 3640
rect 830 3620 850 3630
rect 860 3620 890 3630
rect 990 3620 3020 3630
rect 3080 3620 3140 3630
rect 3210 3620 3270 3630
rect 870 3610 3030 3620
rect 770 3600 780 3610
rect 730 3590 820 3600
rect 850 3590 2940 3610
rect 2950 3600 3030 3610
rect 3090 3610 3150 3620
rect 3210 3610 3310 3620
rect 3390 3610 3430 3630
rect 3500 3620 3660 3630
rect 3680 3620 3690 3630
rect 3500 3610 3690 3620
rect 3717 3620 3770 3630
rect 3810 3621 3830 3630
rect 3850 3621 3900 3640
rect 4060 3630 4490 3640
rect 4540 3630 4560 3640
rect 4670 3630 4740 3660
rect 5270 3650 5290 3660
rect 5310 3660 5400 3670
rect 5410 3660 5480 3670
rect 5310 3650 5460 3660
rect 5490 3650 5550 3670
rect 5640 3660 5730 3690
rect 5830 3680 5890 3690
rect 5940 3680 5960 3690
rect 5830 3670 5910 3680
rect 5930 3670 5970 3680
rect 5830 3660 5970 3670
rect 5630 3650 5730 3660
rect 5860 3650 5990 3660
rect 5260 3630 5300 3650
rect 5310 3640 5470 3650
rect 5310 3630 5480 3640
rect 5490 3630 5510 3650
rect 3810 3620 3900 3621
rect 4050 3620 4530 3630
rect 3717 3610 3780 3620
rect 3820 3610 3910 3620
rect 3090 3600 3160 3610
rect 3250 3600 3320 3610
rect 3390 3600 3440 3610
rect 730 3580 800 3590
rect 840 3580 2940 3590
rect 740 3570 790 3580
rect 830 3570 2940 3580
rect 2970 3590 3040 3600
rect 3090 3590 3190 3600
rect 3260 3590 3320 3600
rect 3400 3590 3440 3600
rect 3490 3590 3810 3610
rect 3822 3609 3910 3610
rect 3830 3600 3910 3609
rect 3820 3590 3920 3600
rect 2970 3580 3050 3590
rect 3090 3580 3100 3590
rect 3120 3580 3200 3590
rect 3270 3580 3330 3590
rect 3420 3580 3430 3590
rect 3480 3580 3920 3590
rect 4060 3590 4560 3620
rect 4690 3610 4740 3630
rect 4850 3610 4860 3630
rect 5250 3610 5510 3630
rect 5540 3640 5560 3650
rect 5620 3640 5720 3650
rect 5870 3640 5990 3650
rect 5540 3620 5568 3640
rect 5616 3630 5710 3640
rect 5530 3618 5568 3620
rect 4600 3600 4610 3610
rect 4690 3600 4720 3610
rect 4600 3590 4620 3600
rect 4690 3590 4700 3600
rect 4750 3590 4770 3610
rect 5260 3600 5430 3610
rect 5460 3600 5470 3610
rect 5530 3600 5570 3618
rect 5580 3610 5600 3615
rect 5620 3610 5710 3630
rect 5870 3630 5970 3640
rect 5870 3620 5910 3630
rect 5880 3610 5910 3620
rect 5940 3620 5970 3630
rect 5940 3610 5950 3620
rect 5580 3600 5690 3610
rect 5260 3590 5420 3600
rect 5540 3590 5690 3600
rect 4060 3580 4570 3590
rect 4600 3580 4630 3590
rect 2970 3570 3100 3580
rect 3140 3570 3210 3580
rect 3270 3570 3340 3580
rect 3470 3570 3930 3580
rect 4060 3570 4370 3580
rect 4380 3570 4620 3580
rect 5260 3570 5430 3590
rect 5550 3580 5690 3590
rect 5550 3570 5700 3580
rect 730 3560 800 3570
rect 810 3560 3090 3570
rect 3150 3560 3210 3570
rect 3280 3560 3350 3570
rect 730 3550 3000 3560
rect 3020 3550 3100 3560
rect 730 3540 2990 3550
rect 3030 3540 3100 3550
rect 3160 3550 3220 3560
rect 3310 3550 3380 3560
rect 3460 3550 3930 3570
rect 4070 3560 4660 3570
rect 5270 3560 5430 3570
rect 4080 3550 4670 3560
rect 5270 3550 5420 3560
rect 5570 3550 5700 3570
rect 5930 3560 5950 3570
rect 6010 3560 6020 3570
rect 5930 3550 5960 3560
rect 5990 3550 6020 3560
rect 3160 3540 3240 3550
rect 3330 3540 3390 3550
rect 3460 3540 3940 3550
rect 4100 3540 4680 3550
rect 4690 3540 4710 3550
rect 5270 3540 5410 3550
rect 750 3530 2990 3540
rect 3040 3530 3110 3540
rect 3160 3530 3170 3540
rect 3190 3530 3260 3540
rect 740 3520 2980 3530
rect 3050 3520 3120 3530
rect 3210 3520 3270 3530
rect 3340 3520 3390 3540
rect 550 3510 560 3520
rect 690 3510 700 3520
rect 730 3510 2970 3520
rect 3070 3510 3150 3520
rect 550 3500 570 3510
rect 720 3500 2980 3510
rect 3090 3500 3160 3510
rect 3220 3500 3280 3520
rect 3350 3510 3410 3520
rect 3380 3500 3420 3510
rect 3450 3500 3940 3540
rect 4110 3530 4710 3540
rect 5280 3530 5410 3540
rect 5600 3530 5700 3550
rect 4120 3520 4420 3530
rect 710 3490 2990 3500
rect 3000 3490 3040 3500
rect 3100 3490 3160 3500
rect 3230 3490 3290 3500
rect 3390 3495 3940 3500
rect 3390 3490 3800 3495
rect 3810 3490 3940 3495
rect 4130 3510 4420 3520
rect 4440 3510 4720 3530
rect 5270 3520 5400 3530
rect 4870 3510 4890 3520
rect 5260 3510 5400 3520
rect 5590 3520 5700 3530
rect 5590 3510 5710 3520
rect 5950 3510 5970 3520
rect 6010 3510 6020 3550
rect 4130 3500 4720 3510
rect 4830 3500 4850 3510
rect 4130 3490 4730 3500
rect 4770 3490 4780 3500
rect 4840 3490 4850 3500
rect 4860 3500 4890 3510
rect 5270 3500 5410 3510
rect 4860 3490 4900 3500
rect 5280 3490 5420 3500
rect 5600 3490 5710 3510
rect 5940 3500 5970 3510
rect 6000 3500 6020 3510
rect 700 3480 3040 3490
rect 3110 3480 3160 3490
rect 3250 3480 3320 3490
rect 3400 3480 3780 3490
rect 3810 3480 3950 3490
rect 4130 3480 4800 3490
rect 4870 3480 4910 3490
rect 5280 3480 5430 3490
rect 5590 3480 5710 3490
rect 690 3470 3050 3480
rect 3110 3470 3170 3480
rect 3280 3470 3330 3480
rect 3410 3470 3770 3480
rect 3810 3470 3960 3480
rect 4130 3470 4490 3480
rect 4510 3470 4800 3480
rect 4890 3470 4910 3480
rect 5250 3470 5400 3480
rect 610 3460 620 3470
rect 680 3460 3050 3470
rect 3120 3460 3210 3470
rect 3280 3460 3340 3470
rect 3410 3460 3970 3470
rect 4130 3460 4810 3470
rect 4890 3460 4980 3470
rect 670 3450 3060 3460
rect 3160 3450 3220 3460
rect 660 3440 3020 3450
rect 3050 3440 3100 3450
rect 3170 3440 3220 3450
rect 3290 3440 3340 3460
rect 3420 3450 3970 3460
rect 4120 3459 4824 3460
rect 4863 3459 4980 3460
rect 3410 3440 3960 3450
rect 4120 3440 4980 3459
rect 610 3420 620 3430
rect 650 3420 3010 3440
rect 3050 3420 3110 3440
rect 3170 3430 3230 3440
rect 3310 3430 3330 3440
rect 3360 3430 3380 3440
rect 3410 3430 3950 3440
rect 4110 3430 4310 3440
rect 4320 3430 4800 3440
rect 250 3410 260 3420
rect 640 3410 3010 3420
rect 3060 3410 3110 3420
rect 3180 3420 3230 3430
rect 3180 3410 3240 3420
rect 3350 3410 3390 3430
rect 3400 3410 3940 3430
rect 4100 3420 4810 3430
rect 4830 3420 4890 3440
rect 4917 3438 4980 3440
rect 4930 3420 4980 3438
rect 5250 3460 5420 3470
rect 5580 3460 5710 3480
rect 5790 3490 5820 3500
rect 5940 3490 6020 3500
rect 5790 3470 5830 3490
rect 5930 3470 6020 3490
rect 5780 3460 5840 3470
rect 5920 3460 6020 3470
rect 5250 3440 5410 3460
rect 5570 3450 5710 3460
rect 5770 3450 5890 3460
rect 5250 3430 5260 3440
rect 5290 3430 5440 3440
rect 5570 3430 5690 3450
rect 5770 3441 5900 3450
rect 4090 3410 4900 3420
rect 630 3400 3020 3410
rect 3070 3408 3110 3410
rect 3070 3400 3099 3408
rect 3220 3400 3280 3410
rect 620 3390 3020 3400
rect 3090 3399 3099 3400
rect 3120 3399 3150 3400
rect 3090 3390 3100 3399
rect 3110 3390 3150 3399
rect 3230 3390 3280 3400
rect 3350 3390 3940 3410
rect 4100 3400 4910 3410
rect 4930 3400 5010 3420
rect 5030 3410 5060 3417
rect 5300 3410 5430 3430
rect 5580 3420 5690 3430
rect 5811 3440 5900 3441
rect 5811 3430 5910 3440
rect 5950 3430 6020 3460
rect 5811 3429 5850 3430
rect 5570 3410 5690 3420
rect 5800 3410 5850 3429
rect 5920 3420 6020 3430
rect 5930 3410 6020 3420
rect 5030 3400 5070 3410
rect 5290 3400 5420 3410
rect 3960 3390 3980 3400
rect 4100 3390 4990 3400
rect 5030 3390 5080 3400
rect 5110 3390 5140 3400
rect 5220 3390 5250 3400
rect 5290 3390 5400 3400
rect 620 3380 3030 3390
rect 3110 3380 3160 3390
rect 3230 3380 3290 3390
rect 610 3360 3040 3380
rect 3110 3370 3170 3380
rect 3240 3370 3290 3380
rect 3120 3360 3170 3370
rect 3250 3360 3290 3370
rect 3370 3370 3990 3390
rect 4110 3380 5000 3390
rect 5020 3380 5080 3390
rect 5120 3380 5170 3390
rect 4110 3370 4940 3380
rect 4970 3370 5090 3380
rect 5130 3370 5190 3380
rect 3370 3360 4000 3370
rect 4120 3360 4950 3370
rect 4980 3360 5230 3370
rect 5310 3360 5400 3390
rect 5560 3370 5690 3410
rect 5810 3400 5830 3410
rect 5940 3390 6020 3410
rect 5930 3380 6020 3390
rect 5940 3370 6020 3380
rect 5560 3360 5680 3370
rect 210 3350 220 3360
rect 600 3350 3050 3360
rect 3120 3350 3189 3360
rect 320 3340 340 3350
rect 590 3340 3050 3350
rect 3130 3340 3190 3350
rect 310 3330 350 3340
rect 590 3330 3060 3340
rect 3156 3339 3220 3340
rect 3170 3330 3220 3339
rect 3300 3333 3340 3360
rect 3370 3350 3960 3360
rect 3970 3350 3990 3360
rect 4130 3350 5050 3360
rect 5060 3350 5230 3360
rect 3360 3333 3480 3350
rect 3490 3340 3910 3350
rect 180 3300 210 3320
rect 230 3310 260 3330
rect 290 3310 350 3330
rect 580 3320 3060 3330
rect 230 3300 250 3310
rect 300 3300 360 3310
rect 130 3290 210 3300
rect 300 3290 350 3300
rect 570 3290 3060 3320
rect 3080 3310 3100 3320
rect 3180 3310 3230 3330
rect 3300 3320 3480 3333
rect 3500 3330 3910 3340
rect 3930 3340 3950 3350
rect 4130 3340 4980 3350
rect 3930 3330 3960 3340
rect 4150 3330 4980 3340
rect 5000 3340 5240 3350
rect 5320 3340 5400 3360
rect 5000 3330 5250 3340
rect 3310 3318 3480 3320
rect 3310 3310 3330 3318
rect 3340 3310 3480 3318
rect 3510 3320 3960 3330
rect 4170 3320 5280 3330
rect 5310 3320 5400 3340
rect 3510 3310 3970 3320
rect 4190 3310 4390 3320
rect 3080 3300 3110 3310
rect 3090 3297 3110 3300
rect 3190 3300 3240 3310
rect 3340 3300 3810 3310
rect 3820 3300 3980 3310
rect 4010 3300 4020 3309
rect 4200 3300 4390 3310
rect 4410 3300 5290 3320
rect 5320 3310 5400 3320
rect 5550 3340 5680 3360
rect 5550 3330 5690 3340
rect 5550 3320 5700 3330
rect 5950 3320 6020 3370
rect 5550 3310 5640 3320
rect 5650 3310 5700 3320
rect 5310 3300 5390 3310
rect 5550 3300 5630 3310
rect 5660 3300 5710 3310
rect 3090 3290 3102 3297
rect 3190 3290 3250 3300
rect 3340 3290 3980 3300
rect 4210 3290 4390 3300
rect 4400 3290 5290 3300
rect 70 3280 110 3290
rect 130 3280 190 3290
rect 280 3280 290 3290
rect 300 3280 340 3290
rect 50 3270 200 3280
rect 210 3270 220 3280
rect 270 3270 290 3280
rect 310 3270 320 3280
rect 560 3270 3070 3290
rect 3230 3280 3280 3290
rect 3340 3280 3990 3290
rect 4010 3280 4020 3290
rect 4220 3280 5290 3290
rect 5330 3280 5390 3300
rect 5540 3290 5607 3300
rect 5650 3290 5710 3300
rect 5970 3290 6020 3320
rect 5540 3280 5590 3290
rect 5620 3280 5630 3288
rect 5650 3280 5720 3290
rect 5980 3280 6020 3290
rect 3240 3270 3290 3280
rect 3340 3270 3500 3280
rect 3520 3270 4020 3280
rect 4230 3270 4420 3280
rect 4450 3270 5300 3280
rect 50 3260 220 3270
rect 280 3260 290 3270
rect 40 3250 220 3260
rect 550 3250 3070 3270
rect 3140 3260 3160 3270
rect 30 3240 80 3250
rect 100 3240 220 3250
rect 540 3240 3080 3250
rect 3130 3240 3170 3260
rect 3250 3250 3290 3270
rect 3330 3260 3500 3270
rect 3530 3260 4020 3270
rect 4240 3260 4410 3270
rect 4450 3260 5310 3270
rect 5340 3260 5370 3280
rect 5380 3260 5390 3280
rect 5550 3270 5580 3280
rect 5620 3270 5730 3280
rect 5800 3270 5810 3280
rect 5990 3270 6020 3280
rect 5630 3260 5740 3270
rect 3320 3250 3500 3260
rect 3260 3240 3290 3250
rect 3310 3240 3510 3250
rect 40 3230 70 3240
rect 110 3230 220 3240
rect 50 3220 190 3230
rect 530 3220 3090 3240
rect 3140 3230 3170 3240
rect 3300 3230 3510 3240
rect 3540 3240 4030 3260
rect 4240 3250 4440 3260
rect 4450 3250 5320 3260
rect 4240 3240 5320 3250
rect 3540 3230 3860 3240
rect 3890 3230 4040 3240
rect 3160 3220 3170 3230
rect 3310 3220 3470 3230
rect 0 3210 190 3220
rect 340 3210 360 3220
rect 530 3210 3100 3220
rect 3410 3210 3470 3220
rect 3490 3220 3860 3230
rect 3900 3220 4040 3230
rect 4250 3230 5320 3240
rect 5340 3250 5390 3260
rect 5340 3240 5400 3250
rect 5410 3240 5420 3250
rect 5570 3240 5580 3260
rect 5660 3250 5740 3260
rect 5790 3250 5810 3270
rect 6000 3250 6020 3270
rect 5660 3240 5710 3250
rect 6010 3240 6020 3250
rect 5340 3230 5420 3240
rect 5670 3230 5710 3240
rect 5810 3230 5820 3240
rect 4250 3220 5420 3230
rect 5490 3220 5500 3230
rect 5640 3220 5650 3230
rect 5660 3220 5720 3230
rect 3490 3210 3820 3220
rect 0 3200 170 3210
rect 340 3200 370 3210
rect 400 3200 430 3210
rect 520 3200 3100 3210
rect 0 3190 130 3200
rect 250 3190 270 3200
rect 0 3180 120 3190
rect 230 3180 260 3190
rect 340 3180 460 3200
rect 480 3190 490 3200
rect 470 3180 500 3190
rect 510 3180 3100 3200
rect 3190 3200 3210 3210
rect 3420 3200 3480 3210
rect 3490 3200 3840 3210
rect 3910 3200 3940 3220
rect 3960 3210 4000 3220
rect 4010 3210 4050 3220
rect 4260 3210 5430 3220
rect 5460 3210 5510 3220
rect 5640 3210 5710 3220
rect 3960 3200 3990 3210
rect 3190 3190 3230 3200
rect 3360 3190 3390 3200
rect 3420 3190 3840 3200
rect 3200 3180 3220 3190
rect 3350 3180 3400 3190
rect 0 3160 110 3180
rect 210 3170 250 3180
rect 330 3170 3110 3180
rect 3280 3170 3300 3180
rect 210 3160 230 3170
rect 300 3160 3110 3170
rect 3270 3160 3300 3170
rect 3350 3170 3410 3180
rect 3420 3170 3520 3190
rect 3550 3180 3840 3190
rect 3860 3190 3870 3200
rect 3920 3190 3940 3200
rect 3970 3190 3990 3200
rect 4010 3200 4040 3210
rect 4120 3200 4130 3210
rect 4010 3190 4030 3200
rect 3860 3180 3880 3190
rect 3920 3180 3950 3190
rect 3960 3180 3990 3190
rect 4260 3180 5360 3210
rect 5370 3200 5530 3210
rect 5640 3200 5700 3210
rect 5380 3190 5530 3200
rect 5630 3190 5690 3200
rect 5380 3180 5540 3190
rect 5630 3180 5700 3190
rect 5810 3180 5820 3190
rect 3350 3160 3400 3170
rect 3430 3162 3520 3170
rect 3560 3170 3890 3180
rect 3920 3170 4000 3180
rect 4210 3170 4220 3180
rect 4260 3170 5530 3180
rect 3430 3160 3531 3162
rect 0 3150 20 3160
rect 0 3130 10 3150
rect 40 3140 130 3160
rect 270 3150 3120 3160
rect 3260 3150 3290 3160
rect 40 3130 160 3140
rect 240 3130 260 3150
rect 280 3130 480 3150
rect 500 3140 3120 3150
rect 3170 3140 3180 3150
rect 490 3130 3130 3140
rect 0 3110 20 3130
rect 40 3120 170 3130
rect 210 3120 220 3130
rect 230 3120 3130 3130
rect 3370 3120 3390 3160
rect 3440 3150 3490 3160
rect 3510 3153 3531 3160
rect 3440 3140 3480 3150
rect 3510 3147 3537 3153
rect 3560 3150 3700 3170
rect 3519 3140 3537 3147
rect 3550 3140 3700 3150
rect 3710 3160 3890 3170
rect 3710 3150 3850 3160
rect 3710 3140 3720 3150
rect 3730 3140 3820 3150
rect 3830 3140 3840 3150
rect 3440 3120 3490 3140
rect 3519 3138 3840 3140
rect 3520 3120 3840 3138
rect 3860 3140 3900 3160
rect 3930 3150 4030 3170
rect 4070 3150 4090 3160
rect 3980 3140 4040 3150
rect 3860 3120 3910 3140
rect 3990 3130 4020 3140
rect 4080 3130 4090 3150
rect 4250 3140 5530 3170
rect 4260 3130 5530 3140
rect 5630 3170 5730 3180
rect 5630 3130 5710 3170
rect 5780 3160 5790 3180
rect 5780 3150 5800 3160
rect 5840 3150 5870 3160
rect 5810 3140 5820 3150
rect 5830 3140 5870 3150
rect 5810 3130 5870 3140
rect 4000 3120 4020 3130
rect 4260 3120 4520 3130
rect 50 3110 190 3120
rect 210 3110 3130 3120
rect 3360 3110 3400 3120
rect 3430 3110 3710 3120
rect 0 3100 10 3110
rect 50 3080 200 3110
rect 210 3100 3140 3110
rect 3360 3100 3410 3110
rect 3420 3100 3710 3110
rect 210 3090 220 3100
rect 240 3090 3140 3100
rect 3280 3090 3310 3100
rect 3360 3090 3540 3100
rect 3560 3090 3710 3100
rect 3720 3110 3810 3120
rect 3820 3110 3850 3120
rect 3720 3100 3850 3110
rect 3860 3110 3920 3120
rect 3860 3100 3930 3110
rect 4000 3100 4030 3120
rect 4260 3110 4480 3120
rect 4490 3110 4520 3120
rect 4530 3120 5530 3130
rect 5600 3120 5710 3130
rect 5820 3120 5880 3130
rect 4530 3110 5520 3120
rect 5610 3110 5710 3120
rect 5840 3110 5880 3120
rect 3720 3090 3960 3100
rect 270 3080 3140 3090
rect 3200 3080 3210 3090
rect 30 3070 180 3080
rect 50 3060 180 3070
rect 270 3070 3150 3080
rect 3190 3070 3220 3080
rect 3280 3070 3320 3090
rect 3360 3080 3530 3090
rect 3360 3070 3410 3080
rect 3430 3070 3530 3080
rect 3560 3070 3960 3090
rect 3990 3070 4040 3100
rect 4080 3080 4090 3090
rect 4260 3080 5520 3110
rect 5630 3090 5700 3110
rect 5840 3100 5870 3110
rect 6010 3100 6020 3110
rect 5850 3090 5870 3100
rect 6000 3090 6020 3100
rect 5640 3080 5700 3090
rect 5840 3080 5870 3090
rect 6010 3080 6020 3090
rect 4080 3070 4100 3080
rect 4270 3070 4520 3080
rect 4530 3070 5520 3080
rect 5670 3070 5700 3080
rect 5830 3070 5870 3080
rect 270 3060 3160 3070
rect 50 3050 190 3060
rect 280 3050 3160 3060
rect 3190 3050 3230 3070
rect 3290 3060 3310 3070
rect 3370 3050 3410 3070
rect 3440 3060 3500 3070
rect 3560 3060 3860 3070
rect 30 3040 190 3050
rect 40 3030 190 3040
rect 290 3040 320 3050
rect 370 3040 3160 3050
rect 3200 3040 3230 3050
rect 290 3030 300 3040
rect 50 3020 90 3030
rect 100 3020 190 3030
rect 380 3020 3160 3040
rect 3210 3020 3230 3040
rect 3380 3040 3410 3050
rect 3450 3040 3500 3060
rect 3550 3050 3860 3060
rect 3520 3040 3860 3050
rect 3870 3040 3950 3070
rect 3990 3060 4030 3070
rect 3380 3030 3420 3040
rect 3450 3030 3950 3040
rect 4000 3050 4030 3060
rect 4280 3050 5510 3070
rect 5680 3060 5690 3070
rect 5820 3060 5870 3070
rect 5670 3050 5690 3060
rect 5830 3050 5870 3060
rect 4000 3040 4020 3050
rect 4290 3040 5520 3050
rect 4000 3030 4010 3040
rect 4290 3030 5530 3040
rect 5650 3030 5680 3050
rect 3380 3020 3430 3030
rect 3450 3020 3960 3030
rect 4300 3020 5530 3030
rect 50 3010 190 3020
rect 40 3003 190 3010
rect 39 3000 190 3003
rect 370 3000 420 3020
rect 430 3000 3170 3020
rect 3210 3010 3240 3020
rect 3380 3010 3860 3020
rect 3880 3010 3960 3020
rect 4160 3010 4170 3020
rect 4300 3010 5540 3020
rect 5860 3010 5870 3050
rect 3210 3000 3250 3010
rect 3380 3000 3450 3010
rect 3460 3000 3860 3010
rect 30 2990 190 3000
rect 390 2990 3180 3000
rect 39 2988 190 2990
rect 50 2980 190 2988
rect 320 2980 360 2990
rect 370 2980 380 2990
rect 50 2970 200 2980
rect 290 2970 380 2980
rect 400 2980 3180 2990
rect 400 2970 3190 2980
rect 3210 2970 3260 3000
rect 3310 2990 3330 3000
rect 3390 2990 3440 3000
rect 3460 2990 3540 3000
rect 3410 2980 3440 2990
rect 3480 2980 3540 2990
rect 3560 2990 3860 3000
rect 3890 2990 3970 3010
rect 4010 3000 4020 3010
rect 4080 3000 4100 3010
rect 4010 2990 4030 3000
rect 4080 2990 4110 3000
rect 4160 2990 4180 3010
rect 4310 3000 5540 3010
rect 4320 2990 5540 3000
rect 3560 2980 3970 2990
rect 4020 2980 4030 2990
rect 4090 2980 4110 2990
rect 4170 2980 4180 2990
rect 3430 2970 3450 2980
rect 3490 2970 3540 2980
rect 3570 2970 3980 2980
rect 4330 2970 5540 2990
rect 50 2960 210 2970
rect 290 2960 300 2970
rect 310 2960 3190 2970
rect 3220 2960 3260 2970
rect 3440 2960 3460 2970
rect 3500 2960 3550 2970
rect 3560 2960 3980 2970
rect 30 2950 210 2960
rect 0 2940 210 2950
rect 330 2940 3190 2960
rect 3230 2950 3260 2960
rect 3450 2950 3480 2960
rect 3500 2950 3980 2960
rect 4340 2960 5470 2970
rect 5510 2960 5540 2970
rect 4340 2950 5480 2960
rect 0 2910 220 2940
rect 290 2930 310 2940
rect 320 2930 3190 2940
rect 3240 2930 3260 2950
rect 3460 2940 3490 2950
rect 3510 2940 3890 2950
rect 3900 2940 3990 2950
rect 3470 2930 3490 2940
rect 240 2919 260 2930
rect 280 2920 3200 2930
rect 280 2919 310 2920
rect 240 2910 310 2919
rect 320 2910 3200 2920
rect 3240 2920 3270 2930
rect 3330 2920 3350 2930
rect 3480 2920 3500 2930
rect 3520 2920 3890 2940
rect 3910 2920 3990 2940
rect 4340 2940 5500 2950
rect 4340 2930 5510 2940
rect 0 2900 210 2910
rect 0 2890 200 2900
rect 0 2880 210 2890
rect 260 2880 3210 2910
rect 3240 2880 3280 2920
rect 3330 2900 3360 2920
rect 3410 2910 3430 2920
rect 3480 2910 3510 2920
rect 3530 2910 3900 2920
rect 3420 2900 3440 2910
rect 3480 2900 3520 2910
rect 3530 2900 3560 2910
rect 3580 2900 3880 2910
rect 3910 2900 4000 2920
rect 4050 2910 4060 2920
rect 4110 2910 4130 2920
rect 4190 2910 4210 2930
rect 4340 2920 5480 2930
rect 5490 2920 5500 2930
rect 4350 2910 5480 2920
rect 4120 2900 4130 2910
rect 3490 2890 3560 2900
rect 3590 2890 4000 2900
rect 4350 2890 5490 2910
rect 5550 2890 5570 2898
rect 3490 2880 3570 2890
rect 3590 2880 4010 2890
rect 0 2870 380 2880
rect 390 2870 3220 2880
rect 3250 2870 3270 2880
rect 3500 2870 3900 2880
rect 3910 2870 4010 2880
rect 4360 2870 5480 2890
rect 0 2860 3220 2870
rect 0 2850 160 2860
rect 180 2850 3220 2860
rect 3510 2860 3900 2870
rect 0 2840 310 2850
rect 330 2840 3230 2850
rect 3360 2840 3380 2850
rect 0 2830 190 2840
rect 210 2830 290 2840
rect 0 2820 200 2830
rect 240 2820 320 2830
rect 340 2820 3230 2840
rect 3270 2830 3290 2840
rect 0 2810 3240 2820
rect 0 2780 270 2810
rect 290 2800 3250 2810
rect 3260 2800 3300 2830
rect 3350 2820 3380 2840
rect 3440 2820 3460 2840
rect 3510 2830 3530 2860
rect 3540 2840 3900 2860
rect 3930 2860 4010 2870
rect 4370 2860 5480 2870
rect 5550 2870 5580 2890
rect 5800 2880 5840 2890
rect 5790 2870 5850 2880
rect 5550 2860 5590 2870
rect 5780 2860 5860 2870
rect 5870 2860 5900 2870
rect 3930 2850 4020 2860
rect 4380 2850 5480 2860
rect 5540 2850 5600 2860
rect 3920 2840 4020 2850
rect 4070 2840 4090 2850
rect 4150 2840 4160 2850
rect 3510 2820 3540 2830
rect 3550 2820 3910 2840
rect 3360 2810 3370 2820
rect 3510 2810 3600 2820
rect 3510 2800 3610 2810
rect 3620 2800 3910 2820
rect 290 2781 300 2800
rect 320 2781 3250 2800
rect 3280 2790 3290 2800
rect 290 2780 3250 2781
rect 0 2770 20 2780
rect 30 2770 280 2780
rect 290 2770 340 2780
rect 360 2770 3250 2780
rect 3520 2780 3910 2800
rect 3930 2810 4030 2840
rect 4070 2830 4100 2840
rect 4220 2830 4240 2850
rect 4390 2840 5480 2850
rect 4410 2830 5480 2840
rect 4080 2820 4090 2830
rect 4420 2810 5480 2830
rect 3930 2790 4040 2810
rect 4430 2800 5480 2810
rect 0 2750 10 2770
rect 30 2760 340 2770
rect 40 2750 290 2760
rect 300 2750 340 2760
rect 350 2750 3260 2770
rect 3380 2760 3400 2770
rect 3290 2750 3310 2760
rect 30 2740 3270 2750
rect 3280 2740 3320 2750
rect 3370 2740 3410 2760
rect 3460 2750 3480 2760
rect 3520 2750 3540 2780
rect 3550 2770 3920 2780
rect 3960 2770 4040 2790
rect 4180 2770 4190 2780
rect 4440 2770 5480 2800
rect 5530 2840 5600 2850
rect 5780 2840 5910 2860
rect 5530 2830 5560 2840
rect 5570 2830 5600 2840
rect 5670 2830 5690 2840
rect 5770 2830 5910 2840
rect 5530 2810 5590 2830
rect 5780 2820 5900 2830
rect 5640 2810 5650 2820
rect 5790 2810 5870 2820
rect 5530 2800 5680 2810
rect 5800 2800 5860 2810
rect 5530 2790 5710 2800
rect 5810 2790 5860 2800
rect 5530 2780 5560 2790
rect 5570 2780 5710 2790
rect 5520 2770 5710 2780
rect 3560 2760 3920 2770
rect 3560 2750 3910 2760
rect 3950 2750 4050 2770
rect 4090 2760 4110 2770
rect 4080 2750 4120 2760
rect 4170 2750 4200 2770
rect 4250 2750 4270 2770
rect 4320 2760 4330 2770
rect 4320 2750 4340 2760
rect 4450 2750 5480 2770
rect 5510 2760 5710 2770
rect 5800 2780 5850 2790
rect 5800 2770 5840 2780
rect 5800 2760 5830 2770
rect 5500 2750 5700 2760
rect 5800 2750 5840 2760
rect 6010 2750 6020 2760
rect 3470 2740 3490 2750
rect 0 2720 290 2740
rect 300 2730 3320 2740
rect 3380 2730 3410 2740
rect 3520 2730 3550 2750
rect 3570 2740 3920 2750
rect 3560 2730 3930 2740
rect 3950 2730 4060 2750
rect 4090 2740 4120 2750
rect 4180 2740 4200 2750
rect 4450 2740 5720 2750
rect 4100 2730 4120 2740
rect 300 2720 330 2730
rect 340 2720 3320 2730
rect 3520 2720 3930 2730
rect 3960 2720 4060 2730
rect 4440 2720 5720 2740
rect 0 2710 40 2720
rect 50 2710 320 2720
rect 340 2710 3290 2720
rect 0 2670 3290 2710
rect 3530 2700 3930 2720
rect 3970 2710 4060 2720
rect 4450 2710 5720 2720
rect 5810 2710 5820 2750
rect 3970 2700 4070 2710
rect 3540 2690 3560 2700
rect 3570 2690 3930 2700
rect 3390 2670 3420 2680
rect 0 2640 3340 2670
rect 3390 2650 3430 2670
rect 3490 2660 3500 2680
rect 3550 2670 3560 2690
rect 3590 2680 3780 2690
rect 3590 2670 3770 2680
rect 3790 2670 3940 2690
rect 3550 2660 3570 2670
rect 3600 2660 3770 2670
rect 3780 2660 3940 2670
rect 3980 2680 4070 2700
rect 4450 2690 5710 2710
rect 4190 2680 4210 2690
rect 4270 2680 4290 2690
rect 4450 2680 4660 2690
rect 4670 2680 5720 2690
rect 5811 2688 5830 2690
rect 3550 2650 3580 2660
rect 3600 2650 3950 2660
rect 3980 2650 4080 2680
rect 4110 2650 4130 2680
rect 4180 2660 4220 2680
rect 4270 2670 4300 2680
rect 4340 2670 4360 2680
rect 4450 2670 5730 2680
rect 5810 2670 5830 2688
rect 6000 2670 6020 2750
rect 4280 2660 4290 2670
rect 4190 2650 4220 2660
rect 3400 2640 3430 2650
rect 3560 2640 3910 2650
rect 3930 2640 3940 2650
rect 3990 2640 4080 2650
rect 0 2630 3330 2640
rect 3570 2630 3590 2640
rect 3620 2630 3780 2640
rect 3790 2630 3950 2640
rect 4000 2630 4080 2640
rect 0 2610 3310 2630
rect 3630 2620 3780 2630
rect 3800 2620 3950 2630
rect 3990 2620 4090 2630
rect 4460 2620 5720 2670
rect 5810 2660 5820 2670
rect 6010 2660 6020 2670
rect 5840 2630 5850 2640
rect 3630 2610 3890 2620
rect 3900 2610 3950 2620
rect 4000 2610 4090 2620
rect 0 2590 3320 2610
rect 3420 2590 3440 2600
rect 0 2580 3350 2590
rect 0 2570 3360 2580
rect 3410 2570 3450 2590
rect 3510 2580 3530 2600
rect 3630 2590 3960 2610
rect 4010 2600 4100 2610
rect 4470 2600 5720 2620
rect 4000 2590 4100 2600
rect 4210 2590 4220 2600
rect 4290 2590 4310 2600
rect 3590 2580 3970 2590
rect 3510 2570 3540 2580
rect 3580 2570 3970 2580
rect 4010 2570 4100 2590
rect 4200 2580 4230 2590
rect 4280 2580 4320 2590
rect 4370 2580 4380 2600
rect 4470 2590 5730 2600
rect 5830 2590 5860 2630
rect 5880 2590 5890 2600
rect 0 2560 80 2570
rect 90 2560 3360 2570
rect 3420 2560 3450 2570
rect 3590 2560 3960 2570
rect 4010 2560 4110 2570
rect 4210 2560 4230 2580
rect 4290 2570 4320 2580
rect 4300 2560 4310 2570
rect 4470 2560 5760 2590
rect 5810 2580 5860 2590
rect 0 2550 3360 2560
rect 3600 2550 3970 2560
rect 0 2530 3350 2550
rect 3610 2540 3620 2550
rect 3630 2540 3970 2550
rect 4020 2540 4110 2560
rect 3630 2530 3980 2540
rect 4040 2530 4110 2540
rect 4470 2540 5570 2560
rect 5580 2550 5770 2560
rect 5580 2540 5780 2550
rect 5820 2540 5860 2580
rect 4470 2530 5560 2540
rect 0 2510 3340 2530
rect 3630 2520 3990 2530
rect 4040 2520 4120 2530
rect 3630 2510 3970 2520
rect 0 2500 3350 2510
rect 0 2410 3380 2500
rect 3430 2490 3470 2510
rect 3530 2490 3550 2510
rect 3600 2500 3620 2510
rect 3630 2500 3980 2510
rect 3440 2470 3470 2490
rect 3540 2480 3550 2490
rect 3590 2490 3980 2500
rect 3590 2480 3990 2490
rect 4040 2480 4130 2520
rect 4480 2510 5560 2530
rect 5580 2530 5850 2540
rect 5580 2520 5840 2530
rect 5590 2510 5830 2520
rect 4180 2490 4190 2510
rect 4240 2480 4250 2500
rect 4300 2480 4330 2510
rect 4390 2500 4400 2510
rect 4390 2490 4410 2500
rect 4400 2480 4410 2490
rect 4480 2490 5550 2510
rect 5590 2500 5610 2510
rect 5630 2500 5840 2510
rect 5590 2490 5620 2500
rect 5630 2490 5810 2500
rect 5820 2490 5860 2500
rect 4480 2480 5560 2490
rect 5590 2480 5870 2490
rect 3600 2460 3990 2480
rect 3630 2450 4000 2460
rect 4050 2450 4130 2480
rect 4310 2470 4320 2480
rect 4480 2470 5570 2480
rect 5590 2470 5900 2480
rect 4490 2460 5610 2470
rect 5630 2460 5910 2470
rect 4500 2450 5600 2460
rect 5630 2450 5907 2460
rect 3630 2440 4010 2450
rect 3640 2430 4020 2440
rect 3460 2410 3490 2420
rect 0 2390 3400 2410
rect 3450 2400 3490 2410
rect 3550 2400 3570 2420
rect 3640 2410 4010 2430
rect 4040 2420 4130 2450
rect 4510 2440 5640 2450
rect 5650 2440 5907 2450
rect 4510 2430 5630 2440
rect 4180 2420 4200 2430
rect 4410 2420 4420 2430
rect 4520 2420 5610 2430
rect 5650 2420 5930 2440
rect 0 2380 3410 2390
rect 3460 2380 3490 2400
rect 3560 2390 3570 2400
rect 3610 2390 4010 2410
rect 4030 2400 4140 2420
rect 4180 2400 4210 2420
rect 4320 2410 4340 2420
rect 4400 2410 4420 2420
rect 4260 2400 4270 2410
rect 4040 2390 4050 2400
rect 3620 2380 4010 2390
rect 4030 2380 4050 2390
rect 4060 2380 4140 2400
rect 4320 2390 4350 2410
rect 4400 2400 4430 2410
rect 4510 2400 5930 2420
rect 4410 2390 4420 2400
rect 4520 2390 5930 2400
rect 4520 2380 5920 2390
rect 0 2340 3400 2380
rect 3620 2370 4140 2380
rect 4530 2370 5920 2380
rect 3630 2360 4140 2370
rect 3640 2350 4150 2360
rect 4540 2350 5910 2370
rect 3650 2340 4150 2350
rect 0 2320 3410 2340
rect 3650 2330 4140 2340
rect 4190 2330 4210 2340
rect 4420 2330 4430 2340
rect 4490 2330 4500 2340
rect 4550 2330 5920 2350
rect 3480 2320 3510 2330
rect 3570 2320 3590 2330
rect 0 2290 3420 2320
rect 3470 2310 3520 2320
rect 3480 2300 3520 2310
rect 3570 2300 3600 2320
rect 3480 2290 3510 2300
rect 3640 2290 4150 2330
rect 4190 2300 4220 2330
rect 4270 2310 4290 2330
rect 4340 2310 4360 2330
rect 4410 2310 4440 2330
rect 4280 2300 4290 2310
rect 4350 2300 4370 2310
rect 4420 2300 4440 2310
rect 4490 2300 4510 2330
rect 4540 2320 5920 2330
rect 4550 2310 5910 2320
rect 4550 2290 5890 2310
rect 0 2240 3430 2290
rect 3650 2280 4160 2290
rect 3650 2270 4150 2280
rect 3660 2260 4150 2270
rect 4560 2270 5900 2290
rect 0 2210 3440 2240
rect 3500 2230 3520 2240
rect 3590 2230 3610 2240
rect 3500 2210 3530 2230
rect 3590 2220 3620 2230
rect 3660 2220 4160 2260
rect 4560 2250 5910 2270
rect 4200 2240 4210 2250
rect 4270 2240 4290 2250
rect 4350 2240 4360 2250
rect 4190 2220 4220 2240
rect 3600 2210 3610 2220
rect 0 2170 3450 2210
rect 3510 2200 3530 2210
rect 3660 2200 4050 2220
rect 4060 2200 4160 2220
rect 4200 2210 4220 2220
rect 4270 2220 4300 2240
rect 4270 2210 4290 2220
rect 4340 2210 4370 2240
rect 4420 2230 4440 2240
rect 4490 2230 4510 2240
rect 4410 2220 4440 2230
rect 4480 2220 4510 2230
rect 4420 2210 4440 2220
rect 4490 2210 4510 2220
rect 4550 2230 4800 2250
rect 4820 2240 5910 2250
rect 4810 2230 5910 2240
rect 4350 2200 4360 2210
rect 4550 2200 5920 2230
rect 3660 2190 4160 2200
rect 4550 2190 4800 2200
rect 4820 2190 5930 2200
rect 3670 2180 4160 2190
rect 4560 2180 4790 2190
rect 4820 2180 5940 2190
rect 3670 2170 4060 2180
rect 0 2150 3460 2170
rect 3670 2160 4050 2170
rect 4070 2160 4170 2180
rect 4550 2170 5950 2180
rect 4550 2160 5970 2170
rect 6010 2160 6020 2170
rect 0 2110 3470 2150
rect 3530 2140 3550 2150
rect 3610 2140 3630 2150
rect 3530 2130 3560 2140
rect 3620 2130 3630 2140
rect 3670 2148 4170 2160
rect 4180 2148 4220 2150
rect 3540 2120 3550 2130
rect 3670 2120 4220 2148
rect 3670 2118 4209 2120
rect 3670 2110 4188 2118
rect 4270 2110 4290 2150
rect 4340 2140 4360 2160
rect 4420 2150 4430 2160
rect 4490 2150 4500 2160
rect 4330 2130 4360 2140
rect 4340 2110 4360 2130
rect 4410 2140 4430 2150
rect 4410 2130 4440 2140
rect 4410 2110 4430 2130
rect 4480 2120 4510 2150
rect 4550 2140 5570 2160
rect 5580 2140 6020 2160
rect 4540 2130 4820 2140
rect 4830 2139 6020 2140
rect 4830 2130 5590 2139
rect 5620 2130 6020 2139
rect 4480 2110 4500 2120
rect 4540 2110 5590 2130
rect 5640 2120 6020 2130
rect 5650 2110 5810 2120
rect 5820 2110 6020 2120
rect 0 2080 3480 2110
rect 3680 2100 4040 2110
rect 4050 2103 4188 2110
rect 4050 2100 4180 2103
rect 3680 2090 4180 2100
rect 0 2050 3490 2080
rect 3550 2060 3570 2070
rect 3690 2060 4180 2090
rect 4550 2100 5600 2110
rect 4550 2070 4600 2100
rect 4610 2070 5600 2100
rect 5640 2090 6020 2110
rect 5640 2080 5800 2090
rect 5810 2080 5830 2090
rect 5840 2080 6020 2090
rect 4540 2060 5600 2070
rect 3540 2050 3570 2060
rect 0 2030 3500 2050
rect 3550 2030 3570 2050
rect 3630 2050 3640 2060
rect 3690 2050 4200 2060
rect 3630 2030 3650 2050
rect 3690 2040 4220 2050
rect 4270 2040 4290 2060
rect 4340 2040 4360 2060
rect 4410 2040 4430 2060
rect 3690 2030 4210 2040
rect 4280 2030 4290 2040
rect 4350 2030 4360 2040
rect 4420 2030 4430 2040
rect 4480 2050 4500 2060
rect 4540 2050 5610 2060
rect 5650 2050 5800 2080
rect 5850 2050 6020 2080
rect 4480 2030 4510 2050
rect 4530 2040 5610 2050
rect 4520 2030 5610 2040
rect 5660 2030 5810 2050
rect 5840 2030 6020 2050
rect 0 2020 3490 2030
rect 3700 2020 4180 2030
rect 4490 2020 4500 2030
rect 4530 2020 5610 2030
rect 0 1990 3500 2020
rect 3700 2010 4190 2020
rect 3710 1990 4190 2010
rect 4540 2000 5610 2020
rect 0 1960 3510 1990
rect 3720 1980 4160 1990
rect 4170 1980 4200 1990
rect 4550 1980 4590 2000
rect 4610 1990 5610 2000
rect 5670 2022 5810 2030
rect 5820 2022 6020 2030
rect 5670 2010 6020 2022
rect 5670 2001 5970 2010
rect 4610 1980 5620 1990
rect 0 1920 3520 1960
rect 3560 1940 3580 1970
rect 3630 1960 3650 1970
rect 3710 1960 4160 1980
rect 4180 1960 4190 1980
rect 3630 1940 3660 1960
rect 3700 1950 4200 1960
rect 3700 1940 3880 1950
rect 3890 1940 3900 1950
rect 3910 1940 4200 1950
rect 4220 1940 4240 1970
rect 4290 1960 4310 1970
rect 4290 1950 4320 1960
rect 4360 1950 4380 1970
rect 4300 1940 4320 1950
rect 4370 1940 4390 1950
rect 4430 1940 4450 1970
rect 4490 1960 4520 1970
rect 4540 1960 5620 1980
rect 4490 1950 5610 1960
rect 5670 1950 5800 2001
rect 5810 2000 5970 2001
rect 5990 2000 6020 2010
rect 5820 1990 5970 2000
rect 6000 1990 6020 2000
rect 5830 1970 5970 1990
rect 5990 1980 6020 1990
rect 5980 1970 6020 1980
rect 5830 1950 6020 1970
rect 4490 1940 4520 1950
rect 3640 1930 3650 1940
rect 3700 1930 4200 1940
rect 4440 1930 4450 1940
rect 4500 1930 4520 1940
rect 4530 1930 5620 1950
rect 5680 1940 5800 1950
rect 5840 1940 6020 1950
rect 5680 1930 6020 1940
rect 0 1900 3530 1920
rect 3710 1910 4210 1930
rect 4500 1920 4510 1930
rect 0 1860 3540 1900
rect 3710 1890 4200 1910
rect 4540 1900 5620 1930
rect 5670 1900 6020 1930
rect 4540 1890 4580 1900
rect 4590 1890 5630 1900
rect 3710 1880 4210 1890
rect 4300 1880 4310 1890
rect 4510 1880 4520 1890
rect 4540 1880 5640 1890
rect 0 1840 3550 1860
rect 3570 1850 3590 1880
rect 3710 1870 4240 1880
rect 3640 1840 3660 1870
rect 3700 1860 4250 1870
rect 3700 1850 4240 1860
rect 4290 1850 4320 1880
rect 4370 1870 4390 1880
rect 4450 1870 4460 1880
rect 4370 1850 4400 1870
rect 4440 1850 4460 1870
rect 4500 1870 5650 1880
rect 4500 1860 5640 1870
rect 5660 1860 6020 1900
rect 4500 1850 6020 1860
rect 3700 1840 4210 1850
rect 4370 1840 4390 1850
rect 0 1810 3560 1840
rect 3710 1830 4210 1840
rect 4510 1830 6020 1850
rect 3720 1820 4220 1830
rect 4520 1820 4530 1830
rect 4550 1820 6020 1830
rect 3750 1810 4220 1820
rect 4550 1810 5710 1820
rect 0 1790 3570 1810
rect 0 1770 3590 1790
rect 3760 1780 4220 1810
rect 4520 1800 4530 1810
rect 4560 1800 5710 1810
rect 5730 1800 6020 1820
rect 4520 1790 4540 1800
rect 4560 1790 6020 1800
rect 0 1760 3600 1770
rect 3650 1760 3660 1780
rect 3720 1770 3740 1780
rect 3750 1770 3880 1780
rect 3890 1770 4250 1780
rect 3710 1760 4250 1770
rect 4300 1760 4320 1790
rect 4370 1780 4390 1790
rect 4450 1780 4470 1790
rect 4370 1760 4400 1780
rect 4440 1760 4470 1780
rect 0 1720 3590 1760
rect 3650 1750 3670 1760
rect 3710 1750 4220 1760
rect 4380 1750 4390 1760
rect 4450 1750 4470 1760
rect 4520 1780 5680 1790
rect 5690 1780 6020 1790
rect 4520 1750 6020 1780
rect 3720 1740 3730 1750
rect 3750 1740 4220 1750
rect 0 1700 3600 1720
rect 3770 1700 4220 1740
rect 4520 1720 4550 1750
rect 4560 1740 6020 1750
rect 4530 1710 4550 1720
rect 4570 1710 6020 1740
rect 0 1670 3610 1700
rect 3660 1680 3670 1690
rect 3770 1680 4230 1700
rect 4390 1690 4400 1700
rect 4460 1690 4470 1700
rect 0 1640 3620 1670
rect 3660 1660 3680 1680
rect 3730 1670 3940 1680
rect 3950 1670 4230 1680
rect 4270 1670 4280 1690
rect 4320 1680 4340 1690
rect 4330 1670 4340 1680
rect 4390 1670 4410 1690
rect 4450 1680 4480 1690
rect 3730 1650 4220 1670
rect 4460 1660 4480 1680
rect 4520 1680 6020 1710
rect 4520 1660 6010 1680
rect 4520 1650 4580 1660
rect 0 1610 3630 1640
rect 3770 1630 4230 1650
rect 3780 1620 4230 1630
rect 4530 1620 4570 1650
rect 4590 1630 6010 1660
rect 0 1590 3640 1610
rect 3780 1600 4240 1620
rect 4530 1610 4580 1620
rect 4590 1610 6020 1630
rect 3740 1590 3750 1600
rect 3770 1590 4240 1600
rect 0 1580 3650 1590
rect 0 1490 3640 1580
rect 3670 1560 3690 1590
rect 3730 1580 3910 1590
rect 3920 1580 4240 1590
rect 4270 1600 4290 1610
rect 4270 1580 4300 1600
rect 4340 1590 4360 1610
rect 4470 1600 4480 1610
rect 4350 1580 4360 1590
rect 4400 1580 4420 1600
rect 3730 1570 3890 1580
rect 3980 1570 4010 1580
rect 4030 1570 4240 1580
rect 4470 1570 4490 1600
rect 4520 1570 6020 1610
rect 3740 1560 3880 1570
rect 4150 1560 4250 1570
rect 4530 1560 6020 1570
rect 3770 1550 3860 1560
rect 3780 1540 3850 1550
rect 3680 1490 3690 1500
rect 3780 1490 3860 1540
rect 4530 1530 4590 1560
rect 4600 1530 6020 1560
rect 4290 1500 4300 1520
rect 4350 1490 4370 1520
rect 4420 1510 4430 1520
rect 4410 1500 4440 1510
rect 4420 1490 4440 1500
rect 0 1480 3650 1490
rect 0 1440 3640 1480
rect 3680 1470 3700 1490
rect 3740 1480 3760 1490
rect 3770 1480 3910 1490
rect 3930 1480 4080 1490
rect 4350 1480 4360 1490
rect 4420 1480 4430 1490
rect 4480 1480 4500 1510
rect 4530 1500 6020 1530
rect 4520 1480 6020 1500
rect 3740 1460 4260 1480
rect 4530 1470 6020 1480
rect 3780 1450 4070 1460
rect 4080 1450 4260 1460
rect 3780 1440 4020 1450
rect 4040 1440 4070 1450
rect 4090 1440 4130 1450
rect 0 1400 3650 1440
rect 3790 1410 4020 1440
rect 4030 1430 4080 1440
rect 4090 1430 4120 1440
rect 4140 1430 4260 1450
rect 4540 1450 6020 1470
rect 4540 1440 4590 1450
rect 4610 1440 6020 1450
rect 4030 1420 4270 1430
rect 4540 1420 6020 1440
rect 4030 1410 4250 1420
rect 4310 1410 4320 1420
rect 3690 1400 3700 1410
rect 0 1320 3660 1400
rect 3680 1380 3700 1400
rect 3750 1400 3770 1410
rect 3790 1400 4250 1410
rect 4370 1400 4380 1420
rect 4430 1410 4440 1420
rect 4430 1400 4450 1410
rect 3750 1390 4130 1400
rect 4140 1390 4270 1400
rect 4430 1390 4440 1400
rect 4490 1390 6020 1420
rect 3750 1380 4250 1390
rect 4500 1380 4520 1390
rect 3750 1370 3760 1380
rect 3790 1350 4270 1380
rect 4540 1370 6020 1390
rect 3800 1330 4280 1350
rect 3800 1320 4270 1330
rect 0 1310 3670 1320
rect 3800 1310 4290 1320
rect 4320 1310 4340 1340
rect 4380 1330 4390 1340
rect 4510 1330 4530 1340
rect 4550 1330 6020 1370
rect 4380 1310 4400 1330
rect 0 1240 3680 1310
rect 3690 1280 3710 1310
rect 3760 1300 4270 1310
rect 4390 1300 4400 1310
rect 4440 1300 4460 1330
rect 3750 1290 4270 1300
rect 4280 1290 4290 1300
rect 4500 1290 6020 1330
rect 3760 1280 4300 1290
rect 3760 1270 4310 1280
rect 3790 1260 4300 1270
rect 3800 1250 4300 1260
rect 4510 1250 4530 1290
rect 3800 1240 4310 1250
rect 4320 1240 4340 1250
rect 4390 1240 4400 1250
rect 4500 1240 4530 1250
rect 4550 1240 6020 1290
rect 0 1220 3690 1240
rect 3800 1220 4340 1240
rect 4380 1220 4400 1240
rect 4450 1230 4460 1240
rect 0 1210 3700 1220
rect 3760 1210 4340 1220
rect 4390 1210 4400 1220
rect 4440 1210 4460 1230
rect 0 1180 3710 1210
rect 3760 1200 4320 1210
rect 4500 1200 6020 1240
rect 3760 1190 4330 1200
rect 0 1150 3700 1180
rect 3770 1170 4330 1190
rect 3810 1160 4330 1170
rect 3810 1150 4090 1160
rect 4110 1150 4330 1160
rect 4500 1150 4530 1200
rect 4540 1190 6020 1200
rect 4550 1150 6020 1190
rect 0 1120 3710 1150
rect 3810 1140 4040 1150
rect 4060 1140 4120 1150
rect 4130 1140 4340 1150
rect 4390 1140 4400 1150
rect 3810 1120 4020 1140
rect 4050 1130 4120 1140
rect 4040 1120 4130 1130
rect 4140 1120 4340 1140
rect 4380 1120 4400 1140
rect 4450 1130 4460 1150
rect 4500 1130 6020 1150
rect 4440 1120 4460 1130
rect 0 1030 3720 1120
rect 3770 1110 4020 1120
rect 3760 1090 4020 1110
rect 4030 1100 4340 1120
rect 4390 1110 4400 1120
rect 4450 1110 4460 1120
rect 4490 1110 6020 1130
rect 4500 1100 6020 1110
rect 4040 1090 4330 1100
rect 3770 1080 4330 1090
rect 3780 1070 3800 1080
rect 3810 1070 4330 1080
rect 4500 1070 4530 1100
rect 4540 1090 6020 1100
rect 3810 1060 4340 1070
rect 4490 1060 4530 1070
rect 4550 1060 6020 1090
rect 3770 1030 3800 1040
rect 3820 1030 4340 1060
rect 4380 1050 4400 1060
rect 4370 1030 4400 1050
rect 0 970 3730 1030
rect 3760 990 4340 1030
rect 4380 1020 4400 1030
rect 4440 1020 4460 1050
rect 4490 1030 6020 1060
rect 4480 1020 6020 1030
rect 3770 980 4340 990
rect 0 940 3740 970
rect 3770 960 3790 980
rect 3780 950 3790 960
rect 3810 950 4340 980
rect 4490 1010 6020 1020
rect 4490 1000 4530 1010
rect 4490 980 4520 1000
rect 4490 970 4530 980
rect 4540 970 6020 1010
rect 4370 960 4390 970
rect 3780 940 3800 950
rect 3810 940 4350 950
rect 0 890 3750 940
rect 3770 930 4350 940
rect 4360 940 4400 960
rect 4440 950 4460 960
rect 4480 950 6020 970
rect 4360 930 4390 940
rect 4440 930 6020 950
rect 3770 910 4340 930
rect 4370 920 4390 930
rect 4450 920 6020 930
rect 4480 910 6020 920
rect 3780 900 4340 910
rect 3790 890 4340 900
rect 0 850 3760 890
rect 3800 880 3810 890
rect 3820 880 4350 890
rect 4490 880 4520 910
rect 4530 880 6020 910
rect 3820 870 4390 880
rect 3830 860 4390 870
rect 3800 850 3810 860
rect 3820 850 4390 860
rect 4440 870 4470 880
rect 4480 870 6020 880
rect 4440 850 6020 870
rect 0 830 3770 850
rect 3790 840 4390 850
rect 3790 830 4380 840
rect 4430 830 6020 850
rect 0 800 4350 830
rect 0 790 3820 800
rect 0 780 1020 790
rect 0 760 1000 780
rect 1040 770 3790 790
rect 3800 780 3820 790
rect 3810 770 3820 780
rect 1040 760 3820 770
rect 3830 790 4350 800
rect 4440 790 4460 830
rect 3830 780 4370 790
rect 4430 780 4460 790
rect 4480 810 6020 830
rect 4480 790 4520 810
rect 4530 790 6020 810
rect 3830 760 4380 780
rect 4430 770 4470 780
rect 4480 770 6020 790
rect 0 750 980 760
rect 1050 750 4380 760
rect 0 740 970 750
rect 1010 740 1020 750
rect 1060 740 4370 750
rect 0 730 960 740
rect 0 720 950 730
rect 1060 720 4350 740
rect 0 700 930 720
rect 1070 710 4350 720
rect 4420 730 6020 770
rect 1070 700 3820 710
rect 3830 700 4360 710
rect 4420 700 4460 730
rect 0 690 920 700
rect 1080 690 3810 700
rect 3840 690 4360 700
rect 4410 690 4460 700
rect 4480 720 6020 730
rect 4480 700 4520 720
rect 4530 700 6020 720
rect 4480 690 6020 700
rect 0 680 910 690
rect 1080 680 3820 690
rect 0 670 890 680
rect 0 660 880 670
rect 1090 660 3820 680
rect 3840 680 4370 690
rect 4400 680 4460 690
rect 4470 680 6020 690
rect 3840 660 4360 680
rect 4400 670 6020 680
rect 4390 660 6020 670
rect 0 650 870 660
rect 1090 650 4360 660
rect 4400 650 6020 660
rect 0 640 860 650
rect 0 630 850 640
rect 1100 630 4350 650
rect 0 620 840 630
rect 0 610 830 620
rect 0 600 820 610
rect 1110 600 4350 630
rect 4400 640 4460 650
rect 4400 600 4450 640
rect 4470 620 6020 650
rect 4480 610 6020 620
rect 0 590 810 600
rect 1120 590 4350 600
rect 4380 590 4450 600
rect 4470 590 6020 610
rect 0 580 800 590
rect 1120 580 4360 590
rect 4370 580 6020 590
rect 0 570 790 580
rect 1120 570 6020 580
rect 0 560 780 570
rect 1130 560 4360 570
rect 4370 560 6020 570
rect 0 550 770 560
rect 1130 550 4350 560
rect 0 540 760 550
rect 1140 540 4350 550
rect 4390 550 6020 560
rect 4390 540 4440 550
rect 4460 540 6020 550
rect 0 530 750 540
rect 0 520 740 530
rect 0 510 730 520
rect 1140 510 4360 540
rect 4400 530 4440 540
rect 4390 510 4440 530
rect 4470 510 6020 540
rect 0 500 720 510
rect 1150 500 4370 510
rect 4380 500 4440 510
rect 4460 500 6020 510
rect 0 490 710 500
rect 0 480 700 490
rect 0 470 690 480
rect 1150 470 6020 500
rect 0 460 680 470
rect 0 450 670 460
rect 0 440 660 450
rect 0 430 650 440
rect 1160 430 4360 470
rect 0 420 640 430
rect 0 410 630 420
rect 1170 410 4360 430
rect 4380 460 6020 470
rect 4380 450 4440 460
rect 4380 420 4430 450
rect 4370 410 4430 420
rect 4460 410 6020 460
rect 0 390 620 410
rect 1170 400 6020 410
rect 0 360 610 390
rect 1180 370 6020 400
rect 1180 360 4430 370
rect 0 340 600 360
rect 0 320 590 340
rect 1190 330 4360 360
rect 4370 330 4420 360
rect 1200 320 4420 330
rect 4450 320 6020 370
rect 0 310 580 320
rect 1200 310 4430 320
rect 4440 310 6020 320
rect 0 290 570 310
rect 1200 300 6020 310
rect 0 270 560 290
rect 1210 280 4970 300
rect 4990 290 6020 300
rect 1210 270 4420 280
rect 4430 270 4970 280
rect 0 260 550 270
rect 0 240 540 260
rect 1210 250 4410 270
rect 0 230 530 240
rect 1220 230 4410 250
rect 4440 230 4970 270
rect 5000 240 6020 290
rect 0 210 520 230
rect 0 200 510 210
rect 0 190 500 200
rect 1220 190 4970 230
rect 0 170 490 190
rect 1230 180 4960 190
rect 1230 170 4410 180
rect 4420 170 4960 180
rect 0 160 480 170
rect 0 150 470 160
rect 0 140 460 150
rect 1230 140 4400 170
rect 4430 150 4960 170
rect 5010 160 6020 240
rect 4420 140 4960 150
rect 0 130 450 140
rect 0 120 430 130
rect 0 110 410 120
rect 1230 110 4960 140
rect 0 100 380 110
rect 0 80 370 100
rect 480 80 500 90
rect 1230 80 4950 110
rect 0 70 380 80
rect 450 70 530 80
rect 0 60 390 70
rect 430 60 560 70
rect 1230 60 4390 80
rect 4410 60 4950 80
rect 0 50 590 60
rect 0 40 640 50
rect 0 30 660 40
rect 1230 30 4940 60
rect 5020 40 6020 160
rect 0 20 700 30
rect 0 10 720 20
rect 0 0 730 10
rect 1240 0 4940 30
rect 5030 0 6020 40
<< end >>
